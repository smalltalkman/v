// Copyright (c) 2026 Alexander Medvednikov. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module transformer

import os
import v2.ast
import v2.pref
import v2.token
import v2.types

// Transformer performs AST-level transformations to simplify
// and normalize code before codegen. This avoids duplicating
// transformation logic across multiple backends (SSA, cleanc, etc.)
pub struct Transformer {
mut:
	pref &pref.Preferences = unsafe { nil }
	env  &types.Environment
	// Current scope for type lookups (walks up scope chain)
	scope &types.Scope = unsafe { nil }
	// Function root scope for registering transformer-created temp variables
	// This allows cleanc to look up temp variable types from the environment
	fn_root_scope &types.Scope = unsafe { nil }
	// Current module for scope lookups
	cur_module string
	// Temp variable counter for desugaring
	temp_counter int
	// Counter for synthesized positions (uses negative values to avoid collision)
	synth_pos_counter int = -1
	// Track needed auto-generated str functions (type_name -> elem_type for arrays)
	needed_str_fns map[string]string
	// Track needed auto-generated array helper functions
	needed_array_contains_fns   map[string]ArrayMethodInfo
	needed_array_index_fns      map[string]ArrayMethodInfo
	needed_array_last_index_fns map[string]ArrayMethodInfo
	// Current function's return type name (for sum type wrapping in returns)
	cur_fn_ret_type_name string
	// When set, match branch values should be wrapped in this sum type
	// (used when a match expression is returned from a function with sum type return)
	sumtype_return_wrap string
	// Smart cast context stack - supports nested smart casts
	smartcast_stack []SmartcastContext
	// Functions that should be elided (conditional compilation, e.g. @[if verbose ?])
	elided_fns map[string]bool
	// Runtime const initializers grouped by module, preserving module discovery order.
	runtime_const_inits_by_mod map[string][]RuntimeConstInit
	runtime_const_modules      []string
	runtime_const_init_fn_name map[string]string
	// Resolved replacement for compile-time pseudo variable @VMODROOT.
	comptime_vmodroot string
	// Statements generated by expression-level expansions (e.g. filter/map)
	// that must be hoisted before the current statement in transform_stmts.
	pending_stmts []ast.Stmt
	// When true, skip lowering value-position IfExpr to temp variable.
	// Set during contexts that already handle IfExpr RHS (e.g. decl_assign).
	skip_if_value_lowering bool
	// For native backends: map interface variable names to their concrete type names.
	// When we see `shape1 := Shape(rect)`, record shape1 → "Rectangle".
	// Used to rewrite interface method calls to direct concrete calls.
	interface_concrete_types map[string]string
}

// SmartcastContext holds info about a single smartcast
struct SmartcastContext {
	expr         string // The expression being smart-cast (e.g., "w.valera")
	variant      string // The variant type name for union member access (e.g., "int", "Kek", "Array_Attribute")
	variant_full string // The full variant name for type casts (e.g., "ast__Kek", "Array_ast__Attribute")
	sumtype      string // The sum type name (e.g., "Valera")
}

struct ArrayMethodInfo {
	array_type string
	elem_type  string
	is_fixed   bool
	fixed_len  int
}

struct RuntimeConstInit {
	name string
	expr ast.Expr
}

pub fn Transformer.new(files []ast.File, env &types.Environment) &Transformer {
	return Transformer.new_with_pref(files, env, unsafe { nil })
}

pub fn Transformer.new_with_pref(files []ast.File, env &types.Environment, p &pref.Preferences) &Transformer {
	mut t := &Transformer{
		pref:                        unsafe { p }
		env:                         unsafe { env }
		needed_str_fns:              map[string]string{}
		needed_array_contains_fns:   map[string]ArrayMethodInfo{}
		needed_array_index_fns:      map[string]ArrayMethodInfo{}
		needed_array_last_index_fns: map[string]ArrayMethodInfo{}
		runtime_const_inits_by_mod:  map[string][]RuntimeConstInit{}
		runtime_const_init_fn_name:  map[string]string{}
	}
	t.comptime_vmodroot = resolve_comptime_vmodroot(files, p)
	return t
}

fn resolve_comptime_vmodroot(files []ast.File, p &pref.Preferences) string {
	if p != unsafe { nil } && p.vroot.len > 0 {
		return p.vroot
	}
	for file in files {
		if root := detect_vmodroot_from_path(file.name) {
			return root
		}
	}
	cwd := os.getwd()
	if root := detect_vmodroot_from_path(cwd) {
		return root
	}
	return ''
}

fn detect_vmodroot_from_path(path string) ?string {
	if path.len == 0 {
		return none
	}
	mut dir := path
	if !os.is_abs_path(dir) {
		cwd := os.getwd()
		if cwd.len > 0 {
			dir = os.join_path(cwd, dir)
		}
	}
	if !os.is_dir(dir) {
		dir = os.dir(dir)
	}
	for _ in 0 .. 16 {
		if os.is_file(os.join_path(dir, 'v.mod')) {
			return dir
		}
		parent := os.dir(dir)
		if parent == dir {
			break
		}
		dir = parent
	}
	return none
}

fn quote_v_string_literal(raw string) string {
	mut escaped := raw.replace('\\', '\\\\')
	escaped = escaped.replace("'", "\\'")
	return "'${escaped}'"
}

fn (t &Transformer) vmodroot_string_literal(pos token.Pos) ast.StringLiteral {
	return ast.StringLiteral{
		kind:  .v
		value: quote_v_string_literal(t.comptime_vmodroot)
		pos:   pos
	}
}

// push_smartcast adds a new smartcast context to the stack
fn (mut t Transformer) push_smartcast(expr string, variant string, sumtype string) {
	t.smartcast_stack << SmartcastContext{
		expr:         expr
		variant:      variant
		variant_full: variant // Default to same as variant
		sumtype:      sumtype
	}
}

// push_smartcast_full adds a smartcast context with separate short and full variant names
fn (mut t Transformer) push_smartcast_full(expr string, variant string, variant_full string, sumtype string) {
	t.smartcast_stack << SmartcastContext{
		expr:         expr
		variant:      variant
		variant_full: variant_full
		sumtype:      sumtype
	}
}

// pop_smartcast removes the most recent smartcast context from the stack
fn (mut t Transformer) pop_smartcast() {
	if t.smartcast_stack.len > 0 {
		t.smartcast_stack = t.smartcast_stack[..t.smartcast_stack.len - 1]
	}
}

// SmartcastRemoveResult holds the removed context and its original index
struct SmartcastRemoveResult {
	ctx SmartcastContext
	idx int
}

// remove_smartcast_for_expr removes the smartcast context for a specific expression
// Returns the removed context or none if not found
fn (mut t Transformer) remove_smartcast_for_expr(expr_str string) ?SmartcastContext {
	if result := t.remove_smartcast_for_expr_with_idx(expr_str) {
		return result.ctx
	}
	return none
}

// remove_smartcast_for_expr_with_idx removes the smartcast context and returns both context and original index
fn (mut t Transformer) remove_smartcast_for_expr_with_idx(expr_str string) ?SmartcastRemoveResult {
	for i := t.smartcast_stack.len - 1; i >= 0; i-- {
		if t.smartcast_stack[i].expr == expr_str {
			ctx := t.smartcast_stack[i]
			// Remove this specific context by creating new slice without this element
			mut new_stack := []SmartcastContext{cap: t.smartcast_stack.len - 1}
			for j, c in t.smartcast_stack {
				if j != i {
					new_stack << c
				}
			}
			t.smartcast_stack = new_stack
			return SmartcastRemoveResult{
				ctx: ctx
				idx: i
			}
		}
	}
	return none
}

// remove_smartcast_ctx_with_idx removes a specific smartcast context and returns
// the removed context with its original index.
fn (mut t Transformer) remove_smartcast_ctx_with_idx(ctx SmartcastContext) ?SmartcastRemoveResult {
	for i := t.smartcast_stack.len - 1; i >= 0; i-- {
		cur := t.smartcast_stack[i]
		if cur.expr == ctx.expr && cur.variant == ctx.variant
			&& cur.variant_full == ctx.variant_full {
			removed := cur
			mut new_stack := []SmartcastContext{cap: t.smartcast_stack.len - 1}
			for j, c in t.smartcast_stack {
				if j != i {
					new_stack << c
				}
			}
			t.smartcast_stack = new_stack
			return SmartcastRemoveResult{
				ctx: removed
				idx: i
			}
		}
	}
	return none
}

// remove_matching_smartcasts temporarily removes all exact copies of ctx.
fn (mut t Transformer) remove_matching_smartcasts(ctx SmartcastContext) []SmartcastRemoveResult {
	mut removed := []SmartcastRemoveResult{}
	for {
		if result := t.remove_smartcast_ctx_with_idx(ctx) {
			removed << result
		} else {
			break
		}
	}
	return removed
}

// restore_smartcasts restores previously removed contexts in original order.
fn (mut t Transformer) restore_smartcasts(removed []SmartcastRemoveResult) {
	for i := removed.len - 1; i >= 0; i-- {
		entry := removed[i]
		t.insert_smartcast_at(entry.idx, entry.ctx)
	}
}

// insert_smartcast_at inserts a smartcast context at a specific position
fn (mut t Transformer) insert_smartcast_at(idx int, ctx SmartcastContext) {
	if idx >= t.smartcast_stack.len {
		// Append at end
		t.smartcast_stack << ctx
	} else {
		// Insert at position
		mut new_stack := []SmartcastContext{cap: t.smartcast_stack.len + 1}
		for i, c in t.smartcast_stack {
			if i == idx {
				new_stack << ctx
			}
			new_stack << c
		}
		// If idx was 0 and loop didn't add, add at beginning
		if idx == 0 && new_stack.len == t.smartcast_stack.len {
			new_stack = [ctx]
			new_stack << t.smartcast_stack
		}
		t.smartcast_stack = new_stack
	}
}

// find_smartcast_for_expr finds the smartcast context that matches the given expression string
// Returns the context or none if not found
fn (t &Transformer) find_smartcast_for_expr(expr_str string) ?SmartcastContext {
	// Empty expression strings are ambiguous (from unhandled AST nodes like IndexExpr)
	// and must never match, as they would incorrectly apply smartcasts to unrelated
	// expressions (e.g., EmptyExpr in enum shorthands like `.assign`).
	if expr_str == '' {
		return none
	}
	// Search from most recent to oldest (reverse order)
	for i := t.smartcast_stack.len - 1; i >= 0; i-- {
		if t.smartcast_stack[i].expr == expr_str {
			return t.smartcast_stack[i]
		}
	}
	return none
}

// has_active_smartcast returns true if there's any active smartcast context
fn (t &Transformer) has_active_smartcast() bool {
	return t.smartcast_stack.len > 0
}

// cur_smartcast_expr returns the current (most recent) smartcast expression or empty string
fn (t &Transformer) cur_smartcast_expr() string {
	if t.smartcast_stack.len > 0 {
		return t.smartcast_stack[t.smartcast_stack.len - 1].expr
	}
	return ''
}

// cur_smartcast_variant returns the current (most recent) smartcast variant or empty string
fn (t &Transformer) cur_smartcast_variant() string {
	if t.smartcast_stack.len > 0 {
		return t.smartcast_stack[t.smartcast_stack.len - 1].variant
	}
	return ''
}

// next_synth_pos returns a unique negative position for synthesized AST nodes
fn (mut t Transformer) next_synth_pos() token.Pos {
	id := t.synth_pos_counter
	t.synth_pos_counter -= 1
	return token.Pos{
		id:     id
		offset: 0
	}
}

// synth_selector creates a typed SelectorExpr with a unique synthesized position
// and registers its type in the environment so downstream passes can resolve it.
fn (mut t Transformer) open_scope() {
	t.scope = types.new_scope(t.scope)
}

// close_scope returns to the parent scope
fn (mut t Transformer) close_scope() {
	if t.scope != unsafe { nil } {
		t.scope = t.scope.parent
	}
}

// is_var_enum checks if a variable's type is an enum
fn (t &Transformer) is_var_enum(name string) ?string {
	typ := t.lookup_var_type(name) or { return none }
	if typ is types.Enum {
		return typ.name
	}
	return none
}

// transform_files transforms all files and returns transformed copies
pub fn (mut t Transformer) transform_files(files []ast.File) []ast.File {
	// Pre-pass: scan all function declarations for conditional compilation attributes
	// to build elided_fns set before transforming call sites
	for file in files {
		for stmt in file.stmts {
			if stmt is ast.FnDecl {
				for attr in stmt.attributes {
					if attr.comptime_cond !is ast.EmptyExpr {
						if !t.eval_comptime_cond(attr.comptime_cond) {
							t.elided_fns[stmt.name] = true
						}
					}
				}
			}
		}
	}
	// Pre-pass: collect const declarations that require runtime initialization.
	t.collect_runtime_const_inits(files)
	mut result := []ast.File{cap: files.len}
	for file in files {
		result << t.transform_file(file)
	}
	t.inject_runtime_const_init_fns(mut result)
	// Generate auto helper functions and add them to the builtin file
	mut generated_fns := []ast.Stmt{}
	if t.needed_str_fns.len > 0 {
		generated_fns << t.generate_str_functions()
	}
	if t.needed_array_contains_fns.len > 0 || t.needed_array_index_fns.len > 0
		|| t.needed_array_last_index_fns.len > 0 {
		generated_fns << t.generate_array_method_functions()
	}
	if generated_fns.len > 0 {
		for i, file in result {
			if file.mod != 'builtin' {
				continue
			}
			mut new_stmts := []ast.Stmt{cap: file.stmts.len}
			for stmt in file.stmts {
				new_stmts << stmt
			}
			for fn_decl in generated_fns {
				new_stmts << fn_decl
			}
			result[i] = ast.File{
				attributes: file.attributes
				mod:        file.mod
				name:       file.name
				stmts:      new_stmts
				imports:    file.imports
			}
			break
		}
	}
	t.inject_main_runtime_const_init_calls(mut result)
	t.propagate_types(result)
	return result
}

fn runtime_const_init_base_name(mod string) string {
	mut suffix := if mod == '' { 'main' } else { mod }
	suffix = suffix.replace('.', '_').replace('-', '_')
	return '__v_init_consts_${suffix}'
}

fn runtime_const_init_call_name(mod string, fn_name string) string {
	if mod != '' && mod != 'main' && mod != 'builtin' {
		return '${mod}__${fn_name}'
	}
	return fn_name
}

fn (mut t Transformer) collect_runtime_const_inits(files []ast.File) {
	for file in files {
		for stmt in file.stmts {
			if stmt is ast.ConstDecl {
				for field in stmt.fields {
					if !t.contains_call_expr(field.value) {
						continue
					}
					if file.mod !in t.runtime_const_inits_by_mod {
						t.runtime_const_modules << file.mod
					}
					mut inits := t.runtime_const_inits_by_mod[file.mod] or { []RuntimeConstInit{} }
					inits << RuntimeConstInit{
						name: field.name
						expr: field.value
					}
					t.runtime_const_inits_by_mod[file.mod] = inits
				}
			}
		}
	}
}

fn (mut t Transformer) transform_expr_in_module(mod string, expr ast.Expr) ast.Expr {
	old_module := t.cur_module
	old_scope := t.scope
	t.cur_module = mod
	if scope := t.get_module_scope(mod) {
		t.scope = scope
	} else {
		t.scope = unsafe { nil }
	}
	transformed := t.transform_expr(expr)
	t.cur_module = old_module
	t.scope = old_scope
	return transformed
}

fn (mut t Transformer) runtime_const_init_fn_stmt(mod string, fn_name string, inits []RuntimeConstInit) ast.Stmt {
	mut stmts := []ast.Stmt{cap: inits.len}
	for item in inits {
		stmts << ast.AssignStmt{
			op:  .assign
			lhs: [ast.Expr(ast.Ident{
				name: item.name
			})]
			rhs: [t.transform_expr_in_module(mod, item.expr)]
		}
	}
	return ast.Stmt(ast.FnDecl{
		name:  fn_name
		typ:   ast.FnType{}
		stmts: stmts
	})
}

fn (mut t Transformer) inject_runtime_const_init_fns(mut files []ast.File) {
	for mod in t.runtime_const_modules {
		inits := t.runtime_const_inits_by_mod[mod] or { []RuntimeConstInit{} }
		if inits.len == 0 {
			continue
		}
		fn_name := runtime_const_init_base_name(mod)
		t.runtime_const_init_fn_name[mod] = fn_name
		fn_stmt := t.runtime_const_init_fn_stmt(mod, fn_name, inits)
		for i, file in files {
			if file.mod != mod {
				continue
			}
			mut new_stmts := []ast.Stmt{cap: file.stmts.len}
			for stmt in file.stmts {
				new_stmts << stmt
			}
			new_stmts << fn_stmt
			files[i] = ast.File{
				attributes: file.attributes
				mod:        file.mod
				name:       file.name
				stmts:      new_stmts
				imports:    file.imports
			}
			break
		}
	}
}

fn (mut t Transformer) inject_main_runtime_const_init_calls(mut files []ast.File) {
	if t.runtime_const_modules.len == 0 {
		return
	}
	mut init_calls := []ast.Stmt{}
	for mod in t.runtime_const_modules {
		fn_name := t.runtime_const_init_fn_name[mod] or { continue }
		call_name := runtime_const_init_call_name(mod, fn_name)
		init_calls << ast.ExprStmt{
			expr: ast.CallExpr{
				lhs: ast.Ident{
					name: call_name
				}
			}
		}
	}
	if init_calls.len == 0 {
		return
	}
	for i, file in files {
		mut changed := false
		mut new_stmts := []ast.Stmt{cap: file.stmts.len}
		for stmt in file.stmts {
			if stmt is ast.FnDecl && !stmt.is_method && stmt.name == 'main' {
				mut fn_stmts := []ast.Stmt{cap: init_calls.len + stmt.stmts.len}
				for call_stmt in init_calls {
					fn_stmts << call_stmt
				}
				for fn_stmt in stmt.stmts {
					fn_stmts << fn_stmt
				}
				new_stmts << ast.FnDecl{
					attributes: stmt.attributes
					is_public:  stmt.is_public
					is_method:  stmt.is_method
					is_static:  stmt.is_static
					receiver:   stmt.receiver
					language:   stmt.language
					name:       stmt.name
					typ:        stmt.typ
					stmts:      fn_stmts
					pos:        stmt.pos
				}
				changed = true
				continue
			}
			new_stmts << stmt
		}
		if changed {
			files[i] = ast.File{
				attributes: file.attributes
				mod:        file.mod
				name:       file.name
				stmts:      new_stmts
				imports:    file.imports
			}
			break
		}
	}
}

fn (mut t Transformer) transform_file(file ast.File) ast.File {
	// Set current module for scope lookups
	t.cur_module = file.mod
	// Set module scope as starting point
	if scope := t.get_module_scope(file.mod) {
		t.scope = scope
	} else {
		t.scope = unsafe { nil }
	}

	mut stmts := []ast.Stmt{cap: file.stmts.len}
	for stmt in file.stmts {
		stmts << t.transform_stmt(stmt)
	}
	return ast.File{
		attributes: file.attributes
		mod:        file.mod
		name:       file.name
		stmts:      stmts
		imports:    file.imports
	}
}

fn (mut t Transformer) transform_stmt(stmt ast.Stmt) ast.Stmt {
	// Check for OrExpr assignment that needs expansion
	if stmt is ast.AssignStmt {
		if expanded := t.try_expand_or_expr_assign(stmt) {
			return expanded
		}
		// Check for map index assignment: m[key] = val -> map__set(&m, &key, &val)
		if transformed := t.try_transform_map_index_assign(stmt) {
			return transformed
		}
	}
	return match stmt {
		ast.AssignStmt {
			t.transform_assign_stmt(stmt)
		}
		ast.BlockStmt {
			ast.BlockStmt{
				stmts: t.transform_stmts(stmt.stmts)
			}
		}
		ast.ComptimeStmt {
			// Unwrap ComptimeStmt - the inner stmt is transformed directly
			t.transform_stmt(stmt.stmt)
		}
		ast.DeferStmt {
			ast.DeferStmt{
				mode:  stmt.mode
				stmts: t.transform_stmts(stmt.stmts)
			}
		}
		ast.ExprStmt {
			// When IfExpr is directly in a statement position (ExprStmt), don't lower
			// to temp variable — it's not used as a value expression.
			is_direct_if := stmt.expr is ast.IfExpr
			saved_skip := t.skip_if_value_lowering
			if is_direct_if {
				t.skip_if_value_lowering = true
			}
			result := ast.Stmt(ast.ExprStmt{
				expr: t.transform_expr(stmt.expr)
			})
			t.skip_if_value_lowering = saved_skip
			result
		}
		ast.FnDecl {
			t.transform_fn_decl(stmt)
		}
		ast.ForStmt {
			t.transform_for_stmt(stmt)
		}
		ast.ForInStmt {
			t.transform_for_in_stmt(stmt)
		}
		ast.ReturnStmt {
			t.transform_return_stmt(stmt)
		}
		ast.ConstDecl {
			t.transform_const_decl(stmt)
		}
		ast.GlobalDecl {
			t.transform_global_decl(stmt)
		}
		ast.AssertStmt {
			ast.AssertStmt{
				expr:  t.transform_expr(stmt.expr)
				extra: stmt.extra
			}
		}
		else {
			stmt
		}
	}
}

fn (mut t Transformer) transform_stmts(stmts []ast.Stmt) []ast.Stmt {
	mut result := []ast.Stmt{cap: stmts.len}
	is_native_be := t.pref != unsafe { nil } && (t.pref.backend == .arm64 || t.pref.backend == .x64)
	for stmt in stmts {
		// Check for OrExpr assignment that expands to multiple statements
		if stmt is ast.AssignStmt {
			// Native backends (arm64/x64): lower interface casts.
			// `shape1 := Shape(rect)` → `shape1 := rect` and record concrete type mapping.
			if is_native_be && stmt.rhs.len == 1 && stmt.lhs.len == 1 && stmt.lhs[0] is ast.Ident
				&& t.is_interface_cast(stmt.rhs[0]) {
				rhs_cast := stmt.rhs[0] as ast.CallOrCastExpr
				lhs_name := (stmt.lhs[0] as ast.Ident).name
				// Get the concrete type name from the value being cast
				if concrete := t.get_expr_type_name(rhs_cast.expr) {
					t.interface_concrete_types[lhs_name] = concrete
				}
				// Replace the interface cast with just the inner value
				result << t.transform_stmt(ast.AssignStmt{
					op:  stmt.op
					lhs: stmt.lhs
					rhs: [rhs_cast.expr]
					pos: stmt.pos
				})
				continue
			}
			if expanded_or_assign := t.try_expand_or_expr_assign_stmts(stmt) {
				// Note: expand_direct_or_expr_assign already transforms expressions internally,
				// so we don't call transform_stmt again to avoid double transformation
				// (which would cause smartcasts to be applied twice)
				result << expanded_or_assign
				continue
			}
			// Check for if-guard expression: x := if r := map[key] { r } else { default }
			if expanded_if_guard_assign := t.try_expand_if_guard_assign_stmts(stmt) {
				for exp_stmt in expanded_if_guard_assign {
					result << t.transform_stmt(exp_stmt)
				}
				continue
			}
			// Check for if-expression assignment: x = if cond { a } else { b }
			// Transform to a statement-form if that assigns in each branch.
			if expanded_if_expr_assign := t.try_expand_if_expr_assign_stmts(stmt) {
				for exp_stmt in expanded_if_expr_assign {
					result << t.transform_stmt(exp_stmt)
				}
				continue
			}
		}
		// Expand compile-time $if at the statement level
		if stmt is ast.ExprStmt {
			if stmt.expr is ast.ComptimeExpr {
				if stmt.expr.expr is ast.IfExpr {
					selected := t.resolve_comptime_if_stmts(stmt.expr.expr)
					// Process through transform_stmts to handle nested $if blocks
					transformed := t.transform_stmts(selected)
					for s in transformed {
						result << s
					}
					continue
				}
			}
		}
		// Check for OrExpr in expression statements (e.g., println(may_fail() or { 0 }))
		if stmt is ast.ExprStmt {
			if expanded_or_stmt := t.try_expand_or_expr_stmt(stmt) {
				// Note: expand_single_or_expr already transforms expressions internally,
				// so we don't call transform_stmt again to avoid double transformation
				// (which would cause interface method _object to be added twice)
				result << expanded_or_stmt
				continue
			}
			// Check for if-guard in expression statements (e.g., if attr := table[name] { ... })
			if expanded_if_guard_stmt := t.try_expand_if_guard_stmt(stmt) {
				// Note: try_expand_if_guard_stmt already transforms expressions internally,
				// so we don't call transform_stmt again to avoid double transformation
				for exp_stmt in expanded_if_guard_stmt {
					result << exp_stmt
				}
				continue
			}
		}
		// Check for flag enum .set() / .clear() calls that need statement-level lowering
		if stmt is ast.ExprStmt {
			if flag_stmt := t.try_transform_flag_enum_set_clear(stmt) {
				result << flag_stmt
				continue
			}
		}
		// Check for OrExpr in return statements
		if stmt is ast.ReturnStmt {
			if expanded_or_return := t.try_expand_or_expr_return(stmt) {
				// Note: expand_single_or_expr already transforms expressions internally,
				// so we don't call transform_stmt again to avoid double transformation.
				// However, transform_expr may have populated pending_stmts (e.g., from
				// lower_if_expr_value), which must be drained before the return stmt.
				if t.pending_stmts.len > 0 {
					// Insert pending_stmts before the last statement (the return).
					for i, es in expanded_or_return {
						if i == expanded_or_return.len - 1 {
							for ps in t.pending_stmts {
								result << ps
							}
							t.pending_stmts.clear()
						}
						result << es
					}
				} else {
					result << expanded_or_return
				}
				continue
			}
			// Check for if-expression in return statements
			// Transform: return if cond { a } else { b }
			// Into: if cond { return a } else { return b }
			if expanded_return_if := t.try_expand_return_if_expr(stmt) {
				for exp_stmt in expanded_return_if {
					result << t.transform_stmt(exp_stmt)
				}
				continue
			}
		}
		// Expand lock/rlock expressions into mutex lock/unlock calls around the body
		if stmt is ast.ExprStmt {
			if stmt.expr is ast.LockExpr {
				result << t.expand_lock_expr(stmt.expr)
				continue
			}
			// Expand map[key] << value to get_and_set + array_push
			if expanded_map_push := t.try_transform_map_index_push(stmt) {
				result << ast.Stmt(expanded_map_push)
				continue
			}
		}
		// Check for map iteration expansion
		if stmt is ast.ForStmt {
			if expanded_for_in_map := t.try_expand_for_in_map(stmt) {
				for exp_stmt in expanded_for_in_map {
					result << t.transform_stmt(exp_stmt)
				}
				continue
			}
		}
		// Transform the statement. Filter/map expression expansions may populate
		// pending_stmts during this call, which must be hoisted before the result.
		result << t.transform_stmt(stmt)
		if t.pending_stmts.len > 0 {
			// Move the just-appended transformed statement to after pending_stmts.
			last := result.pop()
			for ps in t.pending_stmts {
				result << ps
			}
			t.pending_stmts.clear()
			result << last
		}
	}
	return result
}

fn (mut t Transformer) transform_const_decl(decl ast.ConstDecl) ast.ConstDecl {
	mut fields := []ast.FieldInit{cap: decl.fields.len}
	for field in decl.fields {
		fields << ast.FieldInit{
			name:  field.name
			value: t.transform_expr(field.value)
		}
	}
	return ast.ConstDecl{
		is_public: decl.is_public
		fields:    fields
	}
}

fn (mut t Transformer) transform_global_decl(decl ast.GlobalDecl) ast.GlobalDecl {
	mut fields := []ast.FieldDecl{cap: decl.fields.len}
	for field in decl.fields {
		fields << ast.FieldDecl{
			name:       field.name
			typ:        t.transform_expr(field.typ)
			value:      t.transform_expr(field.value)
			attributes: field.attributes
		}
	}
	return ast.GlobalDecl{
		attributes: decl.attributes
		fields:     fields
	}
}

fn (mut t Transformer) transform_assign_stmt(stmt ast.AssignStmt) ast.AssignStmt {
	// Check for string compound assignment: p += x -> p = string__plus(p, x)
	if stmt.op == .plus_assign && stmt.lhs.len == 1 && stmt.rhs.len == 1 {
		lhs_expr := stmt.lhs[0]
		if t.is_string_expr(lhs_expr) {
			// Transform p += x to p = string__plus(p, x)
			return ast.AssignStmt{
				op:  .assign
				lhs: stmt.lhs
				rhs: [
					ast.CallExpr{
						lhs:  ast.Ident{
							name: 'string__plus'
						}
						args: [t.transform_expr(lhs_expr), t.transform_expr(stmt.rhs[0])]
						pos:  stmt.pos
					},
				]
				pos: stmt.pos
			}
		}
	}
	// Lower writes into result/option payload: res.data = v
	if stmt.op == .assign && stmt.lhs.len == 1 && stmt.rhs.len == 1
		&& stmt.lhs[0] is ast.SelectorExpr {
		lhs_sel := stmt.lhs[0] as ast.SelectorExpr
		if lhs_sel.rhs.name == 'data' {
			if lhs_type := t.get_expr_type(lhs_sel.lhs) {
				match lhs_type {
					types.ResultType {
						base_c := t.type_to_c_name(lhs_type.base_type)
						if base_c != '' && base_c != 'void' {
							return ast.AssignStmt{
								op:  .assign
								lhs: [
									t.lower_wrapper_payload_access(t.transform_expr(lhs_sel.lhs),
										base_c),
								]
								rhs: [t.transform_expr(stmt.rhs[0])]
								pos: stmt.pos
							}
						}
					}
					types.OptionType {
						base_c := t.type_to_c_name(lhs_type.base_type)
						if base_c != '' && base_c != 'void' {
							return ast.AssignStmt{
								op:  .assign
								lhs: [
									t.lower_wrapper_payload_access(t.transform_expr(lhs_sel.lhs),
										base_c),
								]
								rhs: [t.transform_expr(stmt.rhs[0])]
								pos: stmt.pos
							}
						}
					}
					else {}
				}
			}
		}
	}

	mut lhs := []ast.Expr{cap: stmt.lhs.len}
	for _, expr in stmt.lhs {
		// For assignment LHS, temporarily remove ALL smartcasts for simple Ident variables.
		// The LHS is the target of the write (the original sum type variable),
		// not the smartcasted variant dereference.
		// Must remove ALL smartcasts (not just one) for nested is-checks on same variable.
		if expr is ast.Ident {
			mut removed_all := []SmartcastRemoveResult{}
			for {
				if removed := t.remove_smartcast_for_expr_with_idx(expr.name) {
					removed_all << removed
				} else {
					break
				}
			}
			lhs << t.transform_expr(expr)
			// Restore in reverse order to maintain original stack positions
			for i := removed_all.len - 1; i >= 0; i-- {
				entry := removed_all[i]
				t.insert_smartcast_at(entry.idx, entry.ctx)
			}
		} else {
			lhs << t.transform_expr(expr)
		}
	}
	is_tuple_lhs := stmt.lhs.len > 1 || (stmt.lhs.len == 1 && stmt.lhs[0] is ast.Tuple)
	// Keep a shallow view of RHS expressions; deep clone can crash on malformed AST payloads.
	mut rhs_src := unsafe { stmt.rhs }
	if is_tuple_lhs && stmt.rhs.len == 1 && stmt.rhs[0] is ast.PostfixExpr {
		postfix := stmt.rhs[0] as ast.PostfixExpr
		if postfix.op in [.not, .question] {
			// For tuple destructuring with `call()!`, keep the raw call expression.
			// Tuple/result unwrapping is handled later by codegen.
			rhs_src = [postfix.expr]
		}
	}
	mut rhs := []ast.Expr{cap: stmt.rhs.len}
	// For decl_assign with IfExpr RHS, skip value-lowering since cleanc
	// already handles this case efficiently (Type name; if (...) { name = a; } else { ... }).
	is_decl_with_if_rhs := stmt.op == .decl_assign && rhs_src.len == 1 && rhs_src[0] is ast.IfExpr
	saved_skip := t.skip_if_value_lowering
	if is_decl_with_if_rhs {
		t.skip_if_value_lowering = true
	}
	for i, expr in rhs_src {
		mut rhs_expr := expr
		// Preserve expected type context for untyped literals like `[]` / `{}` on assignment.
		if i < stmt.lhs.len {
			if lhs_expected := t.get_expr_type(stmt.lhs[i]) {
				rhs_expr = t.resolve_expr_with_expected_type(rhs_expr, lhs_expected)
			} else if stmt.lhs[i] is ast.Ident {
				lhs_name := (stmt.lhs[i] as ast.Ident).name
				lhs_type_name := t.get_var_type_name(lhs_name)
				if lhs_type_name != '' {
					if lhs_expected2 := t.lookup_type(lhs_type_name) {
						rhs_expr = t.resolve_expr_with_expected_type(rhs_expr, lhs_expected2)
					}
				}
			}
		}
		rhs << t.transform_expr(rhs_expr)
	}
	t.skip_if_value_lowering = saved_skip
	// For simple assignments, check if LHS is a sumtype and wrap the RHS if needed
	if stmt.op in [.assign, .decl_assign] && lhs.len == 1 && rhs.len == 1 {
		lhs_name := t.get_var_name(stmt.lhs[0])
		if lhs_name != '' {
			lhs_type_name := t.get_var_type_name(lhs_name)
			if lhs_type_name != '' && t.is_sum_type(lhs_type_name) {
				if wrapped := t.wrap_sumtype_value_transformed(rhs[0], lhs_type_name) {
					rhs = [wrapped]
				}
			}
		}
	}
	return ast.AssignStmt{
		op:  stmt.op
		lhs: lhs
		rhs: rhs
		pos: stmt.pos
	}
}

// get_var_name extracts the variable name from an expression, handling ModifierExpr
fn (t &Transformer) get_var_name(expr ast.Expr) string {
	if expr is ast.Ident {
		return expr.name
	}
	if expr is ast.ModifierExpr {
		// Unwrap modifier (mut, shared, etc.) to get the actual ident
		if expr.expr is ast.Ident {
			return expr.expr.name
		}
	}
	return ''
}

// try_expand_or_expr_assign checks if an assignment has an OrExpr RHS (used by transform_stmt)
// Returns none since expansion is handled by try_expand_or_expr_assign_stmts at the list level
fn (mut t Transformer) try_expand_or_expr_assign(stmt ast.AssignStmt) ?ast.Stmt {
	return none
}

// try_transform_map_index_assign transforms map index assignment to a function call.
// Transforms: m[key] = val -> map__set(&m, &key, &val)
// Also handles compound assignments: m[key] += val -> { tmp = map_get(m,key); tmp += val; map_set(m,key,tmp) }
fn (mut t Transformer) try_transform_map_index_assign(stmt ast.AssignStmt) ?ast.Stmt {
	// Handle compound assignment by converting to: m[key] = m[key] op val
	if stmt.op != .assign && stmt.op != .decl_assign {
		infix_op := match stmt.op {
			.plus_assign { token.Token.plus }
			.minus_assign { token.Token.minus }
			.mul_assign { token.Token.mul }
			.div_assign { token.Token.div }
			.mod_assign { token.Token.mod }
			.and_assign { token.Token.amp }
			.or_assign { token.Token.pipe }
			.xor_assign { token.Token.xor }
			.left_shift_assign { token.Token.left_shift }
			.right_shift_assign { token.Token.right_shift }
			else { return none }
		}
		if stmt.lhs.len != 1 || stmt.rhs.len != 1 {
			return none
		}
		// Convert m[key] op= val to m[key] = m[key] op val
		new_rhs := ast.Expr(ast.InfixExpr{
			lhs: stmt.lhs[0]
			op:  infix_op
			rhs: stmt.rhs[0]
			pos: stmt.pos
		})
		return t.try_transform_map_index_assign(ast.AssignStmt{
			op:  .assign
			lhs: stmt.lhs
			rhs: [new_rhs]
			pos: stmt.pos
		})
	}
	// Check for single LHS that is an IndexExpr
	if stmt.lhs.len != 1 || stmt.rhs.len != 1 {
		return none
	}
	lhs_expr := stmt.lhs[0]
	mut index_expr := ast.IndexExpr{}
	if lhs_expr is ast.IndexExpr {
		index_expr = lhs_expr
	} else if lhs_expr is ast.GenericArgOrIndexExpr {
		// The parser may represent `m[key]` as GenericArgOrIndexExpr due to ambiguity with generic args.
		// For assignment LHS, treat it as an index expression unless lhs is callable (generic specialization).
		if lhs_type := t.get_expr_type(lhs_expr.lhs) {
			if t.is_callable_type(lhs_type) {
				return none
			}
		}
		index_expr = ast.IndexExpr{
			lhs:      lhs_expr.lhs
			expr:     lhs_expr.expr
			is_gated: false
			pos:      lhs_expr.pos
		}
	} else if lhs_expr is ast.GenericArgs {
		// Same ambiguity case: `m[key]` may be parsed as GenericArgs (single arg) rather than IndexExpr.
		if lhs_expr.args.len != 1 {
			return none
		}
		if lhs_type := t.get_expr_type(lhs_expr.lhs) {
			if t.is_callable_type(lhs_type) {
				return none
			}
		}
		index_expr = ast.IndexExpr{
			lhs:      lhs_expr.lhs
			expr:     lhs_expr.args[0]
			is_gated: false
			pos:      lhs_expr.pos
		}
	} else {
		return none
	}
	// Check if the indexed expression is a map and extract key/value types
	map_expr_typ := t.get_expr_type(index_expr.lhs) or { return none }
	map_type := t.unwrap_map_type(map_expr_typ) or { return none }

	// For nested map index assignment (e.g., m['a']['b'] = val), the inner map access
	// must use map__get_and_set to get a pointer to the actual entry, not a copy.
	map_arg := t.map_index_lhs_to_ptr(index_expr.lhs, map_expr_typ)

	// Transform to: { key_tmp := key; val_tmp := val; map__set(&m, &key_tmp, &val_tmp) }
	// Temps are extracted to statement level to avoid scope-escape issues with
	// statement-expression temporaries ({...}) used as function call arguments.
	mut prefix_stmts := []ast.Stmt{}
	key_arg := t.addr_of_with_prefix_temp(index_expr.expr, map_type.key_type, mut prefix_stmts)
	val_arg := t.addr_of_with_prefix_temp(stmt.rhs[0], map_type.value_type, mut prefix_stmts)

	call_stmt := ast.Stmt(ast.ExprStmt{
		expr: ast.CallExpr{
			lhs:  ast.Ident{
				name: 'map__set'
			}
			args: [
				map_arg,
				t.voidptr_cast(key_arg),
				t.voidptr_cast(val_arg),
			]
			pos:  stmt.pos
		}
	})

	if prefix_stmts.len > 0 {
		prefix_stmts << call_stmt
		return ast.BlockStmt{
			stmts: prefix_stmts
		}
	}
	return call_stmt
}

// map_index_lhs_to_ptr generates a pointer expression to a map for use as the first
// argument of map__set. For simple variables (e.g., `m`), it returns `&m`.
// For nested map index expressions (e.g., `outer['key']` where the result is an inner map),
// it uses map__get_and_set to get a pointer to the actual entry in the outer map,
// avoiding the copy-on-read problem that would lose writes to the inner map.
fn (mut t Transformer) map_index_lhs_to_ptr(lhs ast.Expr, lhs_type types.Type) ast.Expr {
	// Check if lhs is a map index expression (nested map case)
	if lhs is ast.IndexExpr {
		outer_type := t.get_expr_type(lhs.lhs) or {
			// Fallback: take address of transformed expression
			return t.addr_of_expr_with_temp(lhs, lhs_type)
		}
		if outer_map := t.unwrap_map_type(outer_type) {
			// Generate: (inner_map_type*) map__get_and_set(&outer, &key, &zero)
			outer_map_arg := t.map_index_lhs_to_ptr(lhs.lhs, outer_type)
			zero_expr := t.zero_value_expr_for_type(outer_map.value_type)
			get_and_set_call := ast.CallExpr{
				lhs:  ast.Ident{
					name: 'map__get_and_set'
				}
				args: [
					outer_map_arg,
					t.voidptr_cast(t.addr_of_expr_with_temp(lhs.expr, outer_map.key_type)),
					t.voidptr_cast(t.addr_of_expr_with_temp(zero_expr, outer_map.value_type)),
				]
			}
			// Cast the voidptr result to the correct map pointer type
			return ast.CastExpr{
				typ:  ast.Ident{
					name: 'map*'
				}
				expr: get_and_set_call
			}
		}
	}
	// Simple case: take address of variable or expression
	if t.is_pointer_type(lhs_type) {
		return t.transform_expr(lhs)
	}
	return t.addr_of_expr_with_temp(lhs, lhs_type)
}

// try_transform_map_index_push transforms map[key] << value to get_and_set + array_push.
// Transforms: m[key] << val -> array__push_noscan((array*)map__get_and_set(&m, &key, &empty), val)
fn (mut t Transformer) try_transform_map_index_push(stmt ast.ExprStmt) ?ast.Stmt {
	if stmt.expr !is ast.InfixExpr {
		return none
	}
	infix := stmt.expr as ast.InfixExpr
	if infix.op != .left_shift {
		return none
	}
	if infix.lhs !is ast.IndexExpr {
		return none
	}
	index_expr := infix.lhs as ast.IndexExpr
	// Check if the indexed expression is a map with array value type
	map_expr_typ := t.get_expr_type(index_expr.lhs) or { return none }
	map_type := t.unwrap_map_type(map_expr_typ) or { return none }
	// Map values can be aliases of arrays (e.g. `[]int` -> `Array_int`). Unwrap aliases.
	mut val_type := map_type.value_type
	for {
		if val_type is types.Alias {
			alias_t := val_type as types.Alias
			val_type = alias_t.base_type
			continue
		}
		break
	}
	if val_type !is types.Array {
		return none
	}
	arr_type := val_type as types.Array
	elem_type_name := t.type_to_c_name(arr_type.elem_type)
	map_arg := if t.is_pointer_type(map_expr_typ) {
		t.transform_expr(index_expr.lhs)
	} else {
		t.addr_of_expr_with_temp(index_expr.lhs, map_expr_typ)
	}
	mut push_exprs := []ast.Expr{cap: 1}
	push_exprs << t.transform_expr(infix.rhs)
	empty_arr := ast.Expr(ast.ArrayInitExpr{
		typ: ast.Expr(ast.Type(ast.ArrayType{
			elem_type: ast.Ident{
				name: elem_type_name
			}
		}))
	})

	// Generate: array__push_noscan(
	//   (array*)map__get_and_set(&m, &key, &empty_array),
	//   (elem_type[1]){value}
	// )
	return ast.ExprStmt{
		expr: ast.CallExpr{
			lhs:  ast.Ident{
				name: 'array__push_noscan'
			}
			args: [
				// (array*)map__get_and_set(&m, &key, &empty_array)
				ast.Expr(ast.CastExpr{
					typ:  ast.Ident{
						name: 'array*'
					}
					expr: ast.CallExpr{
						lhs:  ast.Ident{
							name: 'map__get_and_set'
						}
						args: [
							map_arg,
							// &key
							t.voidptr_cast(t.addr_of_expr_with_temp(index_expr.expr, map_type.key_type)),
							// &empty_array (typed empty array so pushes use the correct element size)
							t.voidptr_cast(t.addr_of_expr_with_temp(empty_arr, map_type.value_type)),
						]
					}
				}),
				// (elem_type[1]){value}
				ast.Expr(ast.ArrayInitExpr{
					typ:   ast.Expr(ast.Type(ast.ArrayType{
						elem_type: ast.Ident{
							name: elem_type_name
						}
					}))
					exprs: push_exprs
				}),
			]
		}
	}
}

// try_expand_or_expr_assign_stmts expands an OrExpr assignment to multiple statements.
// Transforms: a := may_fail(5) or { 0 }
// Into:
//   _t1 := may_fail(5)
//   if _t1.is_error { err := _t1.err; _t1.data = 0 }
//   a := _t1.data
fn (mut t Transformer) try_expand_or_expr_assign_stmts(stmt ast.AssignStmt) ?[]ast.Stmt {
	// Check for assignment with OrExpr somewhere in RHS (single RHS value)
	if stmt.rhs.len != 1 {
		return none
	}
	rhs_expr := stmt.rhs[0]
	// Check if RHS is directly an OrExpr (simple case)
	if rhs_expr is ast.OrExpr {
		return t.expand_direct_or_expr_assign(stmt, rhs_expr)
	}
	// Handle `!` error propagation (PostfixExpr with .not) for native backends.
	// `a := fn()!` expands to: `_t := fn(); if !_t { return 0 }; a := _t`
	// Also handle bare CallExpr/CallOrCastExpr with Result/Option return type
	// (parser sometimes strips PostfixExpr wrapper but the call still needs error propagation)
	if t.pref != unsafe { nil } && (t.pref.backend == .arm64 || t.pref.backend == .x64) {
		mut call_expr := ast.empty_expr
		mut is_error_propagation := false
		if rhs_expr is ast.PostfixExpr {
			postfix := rhs_expr as ast.PostfixExpr
			if postfix.op in [.not, .question] {
				call_expr = postfix.expr
				is_error_propagation = true
			}
		} else if rhs_expr is ast.CallExpr || rhs_expr is ast.CallOrCastExpr {
			// Check if the call returns a Result or Option type
			if ret_type := t.get_expr_type(rhs_expr) {
				if ret_type is types.ResultType || ret_type is types.OptionType {
					call_expr = rhs_expr
					is_error_propagation = true
				}
			}
		}
		if is_error_propagation {
			temp_name := t.gen_temp_name()
			temp_ident := ast.Ident{
				name: temp_name
			}
			mut stmts := []ast.Stmt{}
			// 1. _t := call_expr
			stmts << ast.AssignStmt{
				op:  .decl_assign
				lhs: [ast.Expr(temp_ident)]
				rhs: [t.transform_expr(call_expr)]
				pos: stmt.pos
			}
			// 2. if !_t { return 0 } (error propagation)
			stmts << ast.ExprStmt{
				expr: ast.IfExpr{
					cond:  ast.PrefixExpr{
						op:   .not
						expr: temp_ident
					}
					stmts: [
						ast.Stmt(ast.ReturnStmt{
							exprs: [
								ast.Expr(ast.BasicLiteral{
									value: '0'
									kind:  .number
								}),
							]
						}),
					]
				}
			}
			// 3. a := _t
			stmts << ast.AssignStmt{
				op:  stmt.op
				lhs: stmt.lhs
				rhs: [ast.Expr(temp_ident)]
				pos: stmt.pos
			}
			return stmts
		}
	}
	// Check if RHS contains an OrExpr (nested case like cast(OrExpr))
	if t.expr_has_or_expr(rhs_expr) {
		mut prefix_stmts := []ast.Stmt{}
		new_rhs := t.extract_or_expr(rhs_expr, mut prefix_stmts)
		if prefix_stmts.len == 0 {
			return none
		}
		// Add the final assignment with the extracted expression
		prefix_stmts << ast.AssignStmt{
			op:  stmt.op
			lhs: stmt.lhs
			rhs: [t.transform_expr(new_rhs)]
			pos: stmt.pos
		}
		return prefix_stmts
	}
	return none
}

// expand_direct_or_expr_assign handles the simple case where RHS is directly an OrExpr
fn (mut t Transformer) expand_direct_or_expr_assign(stmt ast.AssignStmt, or_expr ast.OrExpr) ?[]ast.Stmt {
	// The inner expression should be a call that returns Result or Option, OR a map index
	call_expr := or_expr.expr

	// Check for map index with or block: map[key] or { fallback }
	// This is handled specially since it doesn't use Result/Option types
	if call_expr is ast.IndexExpr {
		if map_result := t.try_expand_map_index_or_assign(stmt, or_expr) {
			return map_result
		}
	}

	// Check for string range with or block: s[0..20] or { 'fallback' }
	// The checker types this as `string`, but it needs `string__substr_with_check`
	// which returns `!string` (Result).
	mut is_string_range_or := false
	if call_expr is ast.IndexExpr {
		if call_expr.expr is ast.RangeExpr && t.is_string_expr(call_expr.lhs) {
			is_string_range_or = true
		}
	}

	// Check if expression returns Result or Option using expression-based lookup
	// This works for both function calls and method calls
	mut is_result := t.expr_returns_result(call_expr)
	mut is_option := t.expr_returns_option(call_expr)

	// Fallback to function name lookup for simple function calls
	fn_name := t.get_call_fn_name(call_expr)
	if !is_result && !is_option && fn_name != '' {
		is_result = t.fn_returns_result(fn_name)
		is_option = t.fn_returns_option(fn_name)
	}

	if !is_result && !is_option {
		if is_string_range_or {
			is_result = true
		} else {
			return none
		}
	}

	// Native backends (arm64/x64) don't use Option/Result structs.
	// Expand `a := fn() or { fallback }` to:
	//   _t := fn(); a := if _t { _t } else { fallback }
	if t.pref != unsafe { nil } && (t.pref.backend == .arm64 || t.pref.backend == .x64) {
		temp_name := t.gen_temp_name()
		temp_ident := ast.Ident{
			name: temp_name
		}
		// For ?SumType returns, use _data field check instead of raw truthiness.
		// Sumtypes are {_tag, _data} structs - the first variant has _tag=0,
		// which would be indistinguishable from none (all zeros).
		mut base_type_name := t.get_expr_base_type(call_expr)
		if base_type_name == '' {
			fn_name2 := t.get_call_fn_name(call_expr)
			if fn_name2 != '' {
				base_type_name = t.get_fn_return_base_type(fn_name2)
			}
		}
		is_sumtype_return := base_type_name != '' && t.is_sum_type(base_type_name)
		// Condition expression: _t for simple types, _t._data for sumtypes
		synth_pos2 := t.next_synth_pos()
		cond_expr := if is_sumtype_return {
			t.synth_selector(temp_ident, '_data', types.Type(types.voidptr_))
		} else {
			ast.Expr(temp_ident)
		}
		not_cond_expr := if is_sumtype_return {
			ast.Expr(ast.PrefixExpr{
				op:   .not
				expr: t.synth_selector(ast.Ident{
					name: temp_name
					pos:  synth_pos2
				}, '_data', types.Type(types.voidptr_))
			})
		} else {
			ast.Expr(ast.PrefixExpr{
				op:   .not
				expr: temp_ident
			})
		}
		mut stmts := []ast.Stmt{}
		// 1. _t := call_expr
		stmts << ast.AssignStmt{
			op:  .decl_assign
			lhs: [ast.Expr(temp_ident)]
			rhs: [t.transform_expr(call_expr)]
			pos: stmt.pos
		}
		// 2. Run or-block side effects in else path, then assign
		or_side_effect_stmts, or_value := t.get_or_block_stmts_and_value(or_expr.stmts)
		// If there are side-effect statements (e.g., print_str('error')),
		// wrap them in: if !_t { side_effects... }
		if or_side_effect_stmts.len > 0 {
			stmts << ast.ExprStmt{
				expr: ast.IfExpr{
					cond:  not_cond_expr
					stmts: or_side_effect_stmts
				}
			}
		}
		// 3. a := if _t { _t } else { or_value }
		modified_if := ast.IfExpr{
			cond:      cond_expr
			stmts:     [ast.Stmt(ast.ExprStmt{
				expr: temp_ident
			})]
			else_expr: or_value
		}
		stmts << ast.AssignStmt{
			op:  stmt.op
			lhs: stmt.lhs
			rhs: [ast.Expr(modified_if)]
			pos: stmt.pos
		}
		return stmts
	}

	// Get base type using expression-based lookup first, then fallback
	mut base_type := t.get_expr_base_type(call_expr)
	if base_type == '' && fn_name != '' {
		base_type = t.get_fn_return_base_type(fn_name)
	}
	// String range or-block: the checker typed this as plain string,
	// so base_type lookup fails. Force it to 'string'.
	if is_string_range_or && base_type == '' {
		base_type = 'string'
	}
	is_void_result := base_type == '' || base_type == 'void'
	_ = is_option // suppress unused warning
	// Generate temp variable name
	temp_name := t.gen_temp_name()
	temp_ident := ast.Ident{
		name: temp_name
	}

	// Register temp variable type (the Result/Option wrapper type)
	if wrapper_type := t.get_expr_type(call_expr) {
		if wrapper_type is types.ResultType || wrapper_type is types.OptionType {
			t.register_temp_var(temp_name, wrapper_type)
		}
	} else if ret_type := t.get_method_return_type(call_expr) {
		// Method-call result types are often missing from env expr positions.
		// Register the resolved return wrapper type so cleanc can unwrap `.data`/`.err`.
		if ret_type is types.ResultType || ret_type is types.OptionType {
			t.register_temp_var(temp_name, ret_type)
		}
	} else if fn_name != '' {
		if fn_ret := t.get_fn_return_type(fn_name) {
			if fn_ret is types.ResultType || fn_ret is types.OptionType {
				t.register_temp_var(temp_name, fn_ret)
			}
		}
	}
	// String range or-block: register as _result_string since the checker
	// didn't record a Result type for this expression.
	if is_string_range_or {
		t.register_temp_var(temp_name, types.ResultType{
			base_type: types.string_
		})
	}

	// Build the expanded statements
	mut stmts := []ast.Stmt{}
	// 1. _t1 := call_expr
	transformed_call := t.transform_expr(call_expr)
	// For string range or-blocks, rename string__substr to string__substr_with_check
	// which returns !string (Result) instead of string.
	rhs_expr := if is_string_range_or {
		t.rename_substr_to_checked(transformed_call)
	} else {
		transformed_call
	}
	stmts << ast.AssignStmt{
		op:  .decl_assign
		lhs: [ast.Expr(temp_ident)]
		rhs: [rhs_expr]
		pos: stmt.pos
	}
	// 2. if _t1.is_error { ... } (for Result) or if _t1.state != 0 { ... } (for Option)
	error_cond := if is_result {
		// _t1.is_error
		t.synth_selector(temp_ident, 'is_error', types.Type(types.bool_))
	} else {
		// _t1.state != 0
		ast.Expr(ast.InfixExpr{
			op:  .ne
			lhs: t.synth_selector(temp_ident, 'state', types.Type(types.int_))
			rhs: ast.BasicLiteral{
				kind:  .number
				value: '0'
			}
		})
	}
	// Build the if-block statements
	mut if_stmts := []ast.Stmt{}
	// Keep `err` available in direct-or expansions; some stdlib or-blocks
	// reference it through transformed interpolation paths.
	if_stmts << ast.AssignStmt{
		op:  .decl_assign
		lhs: [ast.Expr(ast.Ident{
			name: 'err'
		})]
		rhs: [
			t.synth_selector(temp_ident, 'err', types.Type(types.Struct{
				name: 'IError'
			})),
		]
	}
	// Check if or-block contains a return statement (control flow)
	if t.or_block_has_return(or_expr.stmts) {
		// Or-block contains return - transform statements here to handle string
		// concatenation and other transformations. This is done here instead of
		// relying on later transform_stmt to avoid double smartcast transformation.
		if_stmts << t.transform_stmts(or_expr.stmts)
	} else if !is_void_result {
		// Or-block provides a value - assign to data (only for non-void results)
		or_side_effect_stmts, or_value := t.get_or_block_stmts_and_value(or_expr.stmts)
		if or_side_effect_stmts.len > 0 {
			if_stmts << or_side_effect_stmts
		}
		// Check if or-value is a void function call (e.g. error_with_pos()).
		// Void calls can't be assigned - treat as control flow instead.
		if t.is_void_call_expr(or_value) {
			if_stmts << ast.ExprStmt{
				expr: or_value
			}
		} else {
			// _t1.data = or_value (the backend will handle proper casting)
			if_stmts << ast.AssignStmt{
				op:  .assign
				lhs: [
					t.synth_selector(temp_ident, 'data', types.Type(types.voidptr_)),
				]
				rhs: [or_value]
			}
		}
	}
	stmts << ast.ExprStmt{
		expr: ast.IfExpr{
			cond:  error_cond
			stmts: if_stmts
		}
	}
	// 3. a := _t1.data (extract value) - only for non-void results
	if !is_void_result {
		// Variable type is already tracked in scope by checker
		stmts << ast.AssignStmt{
			op:  stmt.op
			lhs: stmt.lhs
			rhs: [
				t.synth_selector(temp_ident, 'data', types.Type(types.voidptr_)),
			]
			pos: stmt.pos
		}
	}
	return stmts
}

// gen_temp_name generates a unique temporary variable name
fn (mut t Transformer) gen_temp_name() string {
	t.temp_counter++
	return '_or_t${t.temp_counter}'
}

// register_temp_var registers a temporary variable with its type in fn_root_scope
// This allows cleanc to look up the type from the environment instead of inferring it
fn (mut t Transformer) register_temp_var(name string, typ types.Type) {
	if t.fn_root_scope != unsafe { nil } {
		t.fn_root_scope.insert(name, typ)
	}
}

// gen_filter_temp_name generates a unique temporary variable name for filter expansion
fn (mut t Transformer) gen_filter_temp_name() string {
	t.temp_counter++
	return '_filter_t${t.temp_counter}'
}

// try_expand_filter_or_map_expr expands array.filter(cond) or array.map(body) calls
// in any expression context. Generates temp array + for loop statements, appends them
// to t.pending_stmts, and returns the temp variable ident as the replacement expression.
fn (mut t Transformer) try_expand_filter_or_map_expr(expr ast.Expr) ?ast.Expr {
	method_name, receiver_expr, body_expr := t.get_filter_or_map_call_info(expr) or { return none }
	// Get the array type from the receiver
	array_type := t.get_array_type_str(receiver_expr) or { return none }
	elem_type := array_type['Array_'.len..]
	is_filter := method_name == 'filter'
	// For map, determine result element type from the checker's type info
	mut result_elem := elem_type
	if !is_filter {
		if typ := t.get_expr_type(body_expr) {
			// For function types (fn pointer/literal args), use the return type
			mut resolved_typ := typ
			if typ is types.FnType {
				if rt := typ.get_return_type() {
					resolved_typ = rt
				}
			}
			c_name := t.type_to_c_name(resolved_typ)
			if c_name != '' && c_name != 'void' && c_name != 'int_literal' {
				result_elem = c_name
			}
		}
	}
	// Generate temp variable name
	temp_name := t.gen_filter_temp_name()
	temp_ident := ast.Ident{
		name: temp_name
	}
	it_ident := ast.Ident{
		name: '_filter_it'
	}
	// 1. mut _filter_t1 := []ResultType{cap: 0}
	init_stmt := ast.Stmt(ast.AssignStmt{
		op:  .decl_assign
		lhs: [
			ast.Expr(ast.ModifierExpr{
				kind: .key_mut
				expr: temp_ident
			}),
		]
		rhs: [
			ast.Expr(ast.ArrayInitExpr{
				typ: ast.Expr(ast.Type(ast.ArrayType{
					elem_type: ast.Ident{
						name: result_elem
					}
				}))
				cap: ast.BasicLiteral{
					kind:  .number
					value: '0'
				}
			}),
		]
	})

	// Replace 'it' with '_filter_it' in the body expression.
	// If the body is a function reference (named function), call it with the element:
	// e.g., arr.filter(my_fn) → ... if (my_fn(_filter_it)) { ... }
	// If the body is a FnLiteral/LambdaExpr, inline its body with param replaced:
	// e.g., arr.map(fn (i int) string { return i.str() })
	//   → ... string _v = _filter_it.str(); ...
	transformed_body := if body_expr is ast.Ident && !t.expr_contains_ident_named(body_expr, 'it')
		&& t.is_fn_ident(body_expr) {
		ast.Expr(ast.CallExpr{
			lhs:  t.transform_expr(body_expr)
			args: [ast.Expr(it_ident)]
		})
	} else if body_expr is ast.FnLiteral && body_expr.typ.params.len == 1 {
		// Inline FnLiteral: extract its single return expression and replace param with _filter_it
		// e.g., arr.map(fn (i int) string { return i.str() })
		//   → ... _filter_it.str() ...
		param_name := body_expr.typ.params[0].name
		ret_expr := t.extract_fn_literal_return_expr(body_expr)
		t.replace_named_ident(ret_expr, param_name, '_filter_it')
	} else {
		t.replace_it_ident(body_expr, '_filter_it')
	}

	// Build the for loop body
	mut loop_body := []ast.Stmt{}
	if is_filter {
		// For filter: if cond { array__push(&arr, &it) }
		push_call := ast.CallExpr{
			lhs:  ast.Ident{
				name: 'array__push'
			}
			args: [
				ast.Expr(ast.CastExpr{
					typ:  ast.Ident{
						name: 'array*'
					}
					expr: ast.PrefixExpr{
						op:   .amp
						expr: temp_ident
					}
				}),
				ast.Expr(ast.PrefixExpr{
					op:   .amp
					expr: it_ident
				}),
			]
		}
		loop_body << ast.Stmt(ast.ExprStmt{
			expr: ast.IfExpr{
				cond:  transformed_body
				stmts: [ast.Stmt(ast.ExprStmt{
					expr: push_call
				})]
			}
		})
	} else {
		// For map: mut _filter_v = body; array__push(&arr, &_filter_v)
		t.temp_counter++
		val_name := '_filter_v${t.temp_counter}'
		val_ident := ast.Ident{
			name: val_name
		}
		// mut _filter_v = body_expr
		loop_body << ast.Stmt(ast.AssignStmt{
			op:  .decl_assign
			lhs: [
				ast.Expr(ast.ModifierExpr{
					kind: .key_mut
					expr: val_ident
				}),
			]
			rhs: [ast.Expr(transformed_body)]
		})
		// array__push((array*)&_filter_t, &_filter_v)
		loop_body << ast.Stmt(ast.ExprStmt{
			expr: ast.CallExpr{
				lhs:  ast.Ident{
					name: 'array__push'
				}
				args: [
					ast.Expr(ast.CastExpr{
						typ:  ast.Ident{
							name: 'array*'
						}
						expr: ast.PrefixExpr{
							op:   .amp
							expr: temp_ident
						}
					}),
					ast.Expr(ast.PrefixExpr{
						op:   .amp
						expr: val_ident
					}),
				]
			}
		})
	}

	// 2. for _filter_it in receiver { ... }
	for_stmt := ast.Stmt(ast.ForStmt{
		init:  ast.ForInStmt{
			value: it_ident
			expr:  t.transform_expr(receiver_expr)
		}
		stmts: loop_body
	})

	// Save and restore pending_stmts to prevent transform_stmt(for_stmt) from
	// draining our init_stmt into the for loop body via nested transform_stmts.
	saved_pending := t.pending_stmts.clone()
	t.pending_stmts.clear()
	transformed_init := t.transform_stmt(init_stmt)
	transformed_for := t.transform_stmt(for_stmt)
	t.pending_stmts = saved_pending
	t.pending_stmts << transformed_init
	t.pending_stmts << transformed_for

	// Return the temp variable as the replacement expression
	return temp_ident
}

// get_filter_or_map_call_info extracts info from a filter/map method call.
// Returns (method_name, receiver_expr, body_expr) or none if not a filter/map call.
fn (t &Transformer) get_filter_or_map_call_info(expr ast.Expr) ?(string, ast.Expr, ast.Expr) {
	// Check for CallOrCastExpr: arr.filter(cond) / arr.map(body)
	if expr is ast.CallOrCastExpr {
		if expr.lhs is ast.SelectorExpr {
			sel := expr.lhs as ast.SelectorExpr
			method_name := sel.rhs.name
			if method_name in ['filter', 'map'] {
				return method_name, sel.lhs, expr.expr
			}
		}
	}
	// Check for CallExpr: arr.filter(cond) / arr.map(body)
	if expr is ast.CallExpr {
		if expr.lhs is ast.SelectorExpr {
			sel := expr.lhs as ast.SelectorExpr
			method_name := sel.rhs.name
			if method_name in ['filter', 'map'] && expr.args.len == 1 {
				return method_name, sel.lhs, expr.args[0]
			}
		}
	}
	return none
}

// replace_it_ident replaces all occurrences of 'it' identifier with the given name
fn (t &Transformer) replace_it_ident(expr ast.Expr, new_name string) ast.Expr {
	match expr {
		ast.Ident {
			if expr.name == 'it' {
				return ast.Ident{
					name: new_name
					pos:  expr.pos
				}
			}
			return expr
		}
		ast.InfixExpr {
			return ast.InfixExpr{
				op:  expr.op
				lhs: t.replace_it_ident(expr.lhs, new_name)
				rhs: t.replace_it_ident(expr.rhs, new_name)
				pos: expr.pos
			}
		}
		ast.PrefixExpr {
			return ast.PrefixExpr{
				op:   expr.op
				expr: t.replace_it_ident(expr.expr, new_name)
				pos:  expr.pos
			}
		}
		ast.ParenExpr {
			return ast.ParenExpr{
				expr: t.replace_it_ident(expr.expr, new_name)
				pos:  expr.pos
			}
		}
		ast.CallExpr {
			mut new_args := []ast.Expr{cap: expr.args.len}
			for arg in expr.args {
				new_args << t.replace_it_ident(arg, new_name)
			}
			return ast.CallExpr{
				lhs:  t.replace_it_ident(expr.lhs, new_name)
				args: new_args
				pos:  expr.pos
			}
		}
		ast.CallOrCastExpr {
			return ast.CallOrCastExpr{
				lhs:  t.replace_it_ident(expr.lhs, new_name)
				expr: t.replace_it_ident(expr.expr, new_name)
				pos:  expr.pos
			}
		}
		ast.SelectorExpr {
			return ast.SelectorExpr{
				lhs: t.replace_it_ident(expr.lhs, new_name)
				rhs: expr.rhs
				pos: expr.pos
			}
		}
		ast.IndexExpr {
			return ast.IndexExpr{
				lhs:  t.replace_it_ident(expr.lhs, new_name)
				expr: t.replace_it_ident(expr.expr, new_name)
				pos:  expr.pos
			}
		}
		ast.CastExpr {
			return ast.CastExpr{
				typ:  expr.typ
				expr: t.replace_it_ident(expr.expr, new_name)
				pos:  expr.pos
			}
		}
		ast.StringInterLiteral {
			mut new_inters := []ast.StringInter{cap: expr.inters.len}
			for inter in expr.inters {
				new_inters << ast.StringInter{
					...inter
					expr: t.replace_it_ident(inter.expr, new_name)
				}
			}
			return ast.StringInterLiteral{
				kind:   expr.kind
				values: expr.values
				inters: new_inters
				pos:    expr.pos
			}
		}
		else {
			return expr
		}
	}
}

// replace_named_ident replaces all occurrences of an identifier with the given old_name
// to a new name. This is a generalized version of replace_it_ident.
fn (t &Transformer) replace_named_ident(expr ast.Expr, old_name string, new_name string) ast.Expr {
	match expr {
		ast.Ident {
			if expr.name == old_name {
				return ast.Ident{
					name: new_name
					pos:  expr.pos
				}
			}
			return expr
		}
		ast.InfixExpr {
			return ast.InfixExpr{
				op:  expr.op
				lhs: t.replace_named_ident(expr.lhs, old_name, new_name)
				rhs: t.replace_named_ident(expr.rhs, old_name, new_name)
				pos: expr.pos
			}
		}
		ast.PrefixExpr {
			return ast.PrefixExpr{
				op:   expr.op
				expr: t.replace_named_ident(expr.expr, old_name, new_name)
				pos:  expr.pos
			}
		}
		ast.ParenExpr {
			return ast.ParenExpr{
				expr: t.replace_named_ident(expr.expr, old_name, new_name)
				pos:  expr.pos
			}
		}
		ast.CallExpr {
			mut new_args := []ast.Expr{cap: expr.args.len}
			for arg in expr.args {
				new_args << t.replace_named_ident(arg, old_name, new_name)
			}
			return ast.CallExpr{
				lhs:  t.replace_named_ident(expr.lhs, old_name, new_name)
				args: new_args
				pos:  expr.pos
			}
		}
		ast.CallOrCastExpr {
			return ast.CallOrCastExpr{
				lhs:  t.replace_named_ident(expr.lhs, old_name, new_name)
				expr: t.replace_named_ident(expr.expr, old_name, new_name)
				pos:  expr.pos
			}
		}
		ast.SelectorExpr {
			return ast.SelectorExpr{
				lhs: t.replace_named_ident(expr.lhs, old_name, new_name)
				rhs: expr.rhs
				pos: expr.pos
			}
		}
		ast.IndexExpr {
			return ast.IndexExpr{
				lhs:  t.replace_named_ident(expr.lhs, old_name, new_name)
				expr: t.replace_named_ident(expr.expr, old_name, new_name)
				pos:  expr.pos
			}
		}
		ast.CastExpr {
			return ast.CastExpr{
				typ:  expr.typ
				expr: t.replace_named_ident(expr.expr, old_name, new_name)
				pos:  expr.pos
			}
		}
		ast.StringInterLiteral {
			mut new_inters := []ast.StringInter{cap: expr.inters.len}
			for inter in expr.inters {
				new_inters << ast.StringInter{
					...inter
					expr: t.replace_named_ident(inter.expr, old_name, new_name)
				}
			}
			return ast.StringInterLiteral{
				kind:   expr.kind
				values: expr.values
				inters: new_inters
				pos:    expr.pos
			}
		}
		else {
			return expr
		}
	}
}

// extract_fn_literal_return_expr extracts the single return expression from a FnLiteral.
// For simple FnLiterals like `fn (i int) string { return i.str() }`, extracts `i.str()`.
// Falls back to the body expression of an ExprStmt if no ReturnStmt found.
fn (t &Transformer) extract_fn_literal_return_expr(lit ast.FnLiteral) ast.Expr {
	for stmt in lit.stmts {
		if stmt is ast.ReturnStmt {
			if stmt.exprs.len > 0 {
				return stmt.exprs[0]
			}
		}
		// Also handle expression statements (implicit return)
		if stmt is ast.ExprStmt {
			return stmt.expr
		}
	}
	// Fallback: return a zero literal (should not be reached for valid FnLiterals)
	return ast.BasicLiteral{
		kind:  .number
		value: '0'
	}
}

// or_block_has_return checks if the or-block contains a control flow statement
// (return, continue, break, panic, exit)
fn (t &Transformer) or_block_has_return(stmts []ast.Stmt) bool {
	for stmt in stmts {
		if stmt is ast.ReturnStmt {
			return true
		}
		if stmt is ast.FlowControlStmt {
			// break, continue, goto
			return true
		}
		if stmt is ast.ExprStmt {
			// Check for panic() or exit() calls
			if stmt.expr is ast.CallExpr {
				if stmt.expr.lhs is ast.Ident {
					name := stmt.expr.lhs.name
					if name in ['panic', 'exit'] {
						return true
					}
				}
			} else if stmt.expr is ast.CallOrCastExpr {
				if stmt.expr.lhs is ast.Ident {
					name := stmt.expr.lhs.name
					if name in ['panic', 'exit'] {
						return true
					}
				}
			}
			// Check for nested OrExpr that contains control flow
			// e.g., scopes[k1] or { scopes[k2] or { return -999 } }
			if stmt.expr is ast.OrExpr {
				or_expr := stmt.expr as ast.OrExpr
				if t.or_block_has_return(or_expr.stmts) {
					return true
				}
			}
		}
	}
	return false
}

fn (t &Transformer) stmt_uses_ident(stmt ast.Stmt, name string) bool {
	match stmt {
		ast.AssignStmt {
			for lhs in stmt.lhs {
				if t.expr_contains_ident_named(lhs, name) {
					return true
				}
			}
			for rhs in stmt.rhs {
				if t.expr_contains_ident_named(rhs, name) {
					return true
				}
			}
		}
		ast.ExprStmt {
			return t.expr_contains_ident_named(stmt.expr, name)
		}
		ast.ReturnStmt {
			for expr in stmt.exprs {
				if t.expr_contains_ident_named(expr, name) {
					return true
				}
			}
		}
		ast.ForStmt {
			if t.stmt_uses_ident(stmt.init, name) || t.expr_contains_ident_named(stmt.cond, name)
				|| t.stmt_uses_ident(stmt.post, name) {
				return true
			}
			for body_stmt in stmt.stmts {
				if t.stmt_uses_ident(body_stmt, name) {
					return true
				}
			}
		}
		ast.BlockStmt {
			for body_stmt in stmt.stmts {
				if t.stmt_uses_ident(body_stmt, name) {
					return true
				}
			}
		}
		ast.DeferStmt {
			for body_stmt in stmt.stmts {
				if t.stmt_uses_ident(body_stmt, name) {
					return true
				}
			}
		}
		else {}
	}
	return false
}

fn (t &Transformer) stmts_use_ident(stmts []ast.Stmt, name string) bool {
	for stmt in stmts {
		if t.stmt_uses_ident(stmt, name) {
			return true
		}
	}
	return false
}

// get_or_block_value extracts the value expression from an or-block
// The value is typically the last expression statement, or 0/default for empty blocks
fn (mut t Transformer) get_or_block_value(stmts []ast.Stmt) ast.Expr {
	_, value := t.get_or_block_stmts_and_value(stmts)
	return value
}

// get_or_block_stmts_and_value extracts side-effect statements and fallback value
// from an or-block. Side effects are all statements before the trailing value expr.
fn (mut t Transformer) get_or_block_stmts_and_value(stmts []ast.Stmt) ([]ast.Stmt, ast.Expr) {
	if stmts.len == 0 {
		return []ast.Stmt{}, ast.Expr(ast.BasicLiteral{
			kind:  .number
			value: '0'
		})
	}
	last := stmts[stmts.len - 1]
	if last is ast.ExprStmt {
		side_effects := if stmts.len > 1 {
			t.transform_stmts(stmts[..stmts.len - 1])
		} else {
			[]ast.Stmt{}
		}
		return side_effects, t.transform_expr(last.expr)
	}
	return t.transform_stmts(stmts), ast.Expr(ast.BasicLiteral{
		kind:  .number
		value: '0'
	})
}

// try_expand_or_expr_stmt handles OrExpr in expression statements like println(may_fail() or { 0 })
// Transforms: println(may_fail(5) or { 0 })
// Into:
//   _t1 := may_fail(5)
//   if _t1.is_error { err := _t1.err; _t1.data = 0 }
//   println(_t1.data)
fn (mut t Transformer) try_expand_or_expr_stmt(stmt ast.ExprStmt) ?[]ast.Stmt {
	// Check if expression contains any OrExpr
	if !t.expr_has_or_expr(stmt.expr) {
		return none
	}
	// Extract OrExpr and get prefix statements + transformed expression
	mut prefix_stmts := []ast.Stmt{}
	new_expr := t.extract_or_expr(stmt.expr, mut prefix_stmts)
	if prefix_stmts.len == 0 {
		return none
	}
	// Add the final expression statement
	prefix_stmts << ast.ExprStmt{
		expr: t.transform_expr(new_expr)
	}
	return prefix_stmts
}

// try_expand_or_expr_return handles OrExpr in return statements
// Transforms: return may_fail(5) or { 0 }
// Into:
//   _t1 := may_fail(5)
//   if _t1.is_error { err := _t1.err; _t1.data = 0 }
//   return _t1.data
fn (mut t Transformer) try_expand_or_expr_return(stmt ast.ReturnStmt) ?[]ast.Stmt {
	// Check if any return expression contains OrExpr
	mut has_or_expr := false
	for expr in stmt.exprs {
		if t.expr_has_or_expr(expr) {
			has_or_expr = true
			break
		}
	}
	if !has_or_expr {
		return none
	}
	// Extract OrExpr from all return expressions
	mut prefix_stmts := []ast.Stmt{}
	mut new_exprs := []ast.Expr{cap: stmt.exprs.len}
	for expr in stmt.exprs {
		new_expr := t.extract_or_expr(expr, mut prefix_stmts)
		new_exprs << t.transform_expr(new_expr)
	}
	if prefix_stmts.len == 0 {
		return none
	}
	// Add the final return statement
	prefix_stmts << ast.ReturnStmt{
		exprs: new_exprs
	}
	return prefix_stmts
}

// expr_has_or_expr checks if an expression contains any OrExpr
fn (t &Transformer) expr_has_or_expr(expr ast.Expr) bool {
	if expr is ast.OrExpr {
		return true
	}
	match expr {
		ast.CallExpr {
			for arg in expr.args {
				if t.expr_has_or_expr(arg) {
					return true
				}
			}
		}
		ast.CallOrCastExpr {
			if t.expr_has_or_expr(expr.expr) {
				return true
			}
		}
		ast.InfixExpr {
			if t.expr_has_or_expr(expr.lhs) || t.expr_has_or_expr(expr.rhs) {
				return true
			}
		}
		ast.PrefixExpr {
			if t.expr_has_or_expr(expr.expr) {
				return true
			}
		}
		ast.ParenExpr {
			if t.expr_has_or_expr(expr.expr) {
				return true
			}
		}
		ast.IndexExpr {
			if t.expr_has_or_expr(expr.lhs) || t.expr_has_or_expr(expr.expr) {
				return true
			}
		}
		ast.SelectorExpr {
			if t.expr_has_or_expr(expr.lhs) {
				return true
			}
		}
		ast.CastExpr {
			if t.expr_has_or_expr(expr.expr) {
				return true
			}
		}
		ast.IfExpr {
			if t.expr_has_or_expr(expr.cond) {
				return true
			}
			if t.expr_has_or_expr(expr.else_expr) {
				return true
			}
			// Note: stmts inside IfExpr are handled separately by transform_stmts
		}
		ast.MatchExpr {
			if t.expr_has_or_expr(expr.expr) {
				return true
			}
		}
		ast.ArrayInitExpr {
			for e in expr.exprs {
				if t.expr_has_or_expr(e) {
					return true
				}
			}
		}
		ast.InitExpr {
			for field in expr.fields {
				if t.expr_has_or_expr(field.value) {
					return true
				}
			}
		}
		else {}
	}
	return false
}

// extract_or_expr extracts OrExpr from an expression tree.
// It generates prefix statements for the OrExpr expansion and returns the expression
// with OrExpr replaced by the temp variable's data access.
fn (mut t Transformer) extract_or_expr(expr ast.Expr, mut prefix_stmts []ast.Stmt) ast.Expr {
	// If this is an OrExpr, expand it directly
	if expr is ast.OrExpr {
		return t.expand_single_or_expr(expr, mut prefix_stmts)
	}
	// Recursively check sub-expressions
	match expr {
		ast.CallExpr {
			mut new_args := []ast.Expr{cap: expr.args.len}
			for arg in expr.args {
				new_args << t.extract_or_expr(arg, mut prefix_stmts)
			}
			return ast.CallExpr{
				lhs:  expr.lhs
				args: new_args
				pos:  expr.pos
			}
		}
		ast.CallOrCastExpr {
			new_inner := t.extract_or_expr(expr.expr, mut prefix_stmts)
			return ast.CallOrCastExpr{
				lhs:  expr.lhs
				expr: new_inner
				pos:  expr.pos
			}
		}
		ast.InfixExpr {
			new_lhs := t.extract_or_expr(expr.lhs, mut prefix_stmts)
			new_rhs := t.extract_or_expr(expr.rhs, mut prefix_stmts)
			return ast.InfixExpr{
				op:  expr.op
				lhs: new_lhs
				rhs: new_rhs
				pos: expr.pos
			}
		}
		ast.PrefixExpr {
			new_inner := t.extract_or_expr(expr.expr, mut prefix_stmts)
			return ast.PrefixExpr{
				op:   expr.op
				expr: new_inner
				pos:  expr.pos
			}
		}
		ast.ParenExpr {
			new_inner := t.extract_or_expr(expr.expr, mut prefix_stmts)
			return ast.ParenExpr{
				expr: new_inner
				pos:  expr.pos
			}
		}
		ast.IndexExpr {
			new_lhs := t.extract_or_expr(expr.lhs, mut prefix_stmts)
			new_idx := t.extract_or_expr(expr.expr, mut prefix_stmts)
			return ast.IndexExpr{
				lhs:      new_lhs
				expr:     new_idx
				is_gated: expr.is_gated
			}
		}
		ast.SelectorExpr {
			new_lhs := t.extract_or_expr(expr.lhs, mut prefix_stmts)
			return ast.SelectorExpr{
				lhs: new_lhs
				rhs: expr.rhs
				pos: expr.pos
			}
		}
		ast.CastExpr {
			new_inner := t.extract_or_expr(expr.expr, mut prefix_stmts)
			return ast.CastExpr{
				typ:  expr.typ
				expr: new_inner
				pos:  expr.pos
			}
		}
		ast.IfExpr {
			new_cond := t.extract_or_expr(expr.cond, mut prefix_stmts)
			new_else := t.extract_or_expr(expr.else_expr, mut prefix_stmts)
			return ast.IfExpr{
				cond:      new_cond
				stmts:     expr.stmts // stmts are processed separately by transform_stmts
				else_expr: new_else
				pos:       expr.pos
			}
		}
		ast.MatchExpr {
			new_matched := t.extract_or_expr(expr.expr, mut prefix_stmts)
			return ast.MatchExpr{
				expr:     new_matched
				branches: expr.branches
				pos:      expr.pos
			}
		}
		ast.ArrayInitExpr {
			mut new_exprs := []ast.Expr{cap: expr.exprs.len}
			for e in expr.exprs {
				new_exprs << t.extract_or_expr(e, mut prefix_stmts)
			}
			return ast.ArrayInitExpr{
				typ:   expr.typ
				exprs: new_exprs
			}
		}
		ast.InitExpr {
			mut new_fields := []ast.FieldInit{cap: expr.fields.len}
			for field in expr.fields {
				new_fields << ast.FieldInit{
					name:  field.name
					value: t.extract_or_expr(field.value, mut prefix_stmts)
				}
			}
			return ast.InitExpr{
				typ:    expr.typ
				fields: new_fields
			}
		}
		else {
			return expr
		}
	}
}

// expand_single_or_expr expands a single OrExpr and returns the data access expression
fn (mut t Transformer) expand_single_or_expr(or_expr ast.OrExpr, mut prefix_stmts []ast.Stmt) ast.Expr {
	call_expr := or_expr.expr

	// Check for map index with or block: map[key] or { fallback }
	if result := t.try_expand_map_index_or(or_expr, mut prefix_stmts) {
		return result
	}

	// Check for string range with or block: s[0..20] or { 'fallback' }
	mut is_string_range_or := false
	if call_expr is ast.IndexExpr {
		if call_expr.expr is ast.RangeExpr && t.is_string_expr(call_expr.lhs) {
			is_string_range_or = true
		}
	}

	// Check if expression returns Result or Option using expression-based lookup
	// This works for both function calls and method calls
	mut is_result := t.expr_returns_result(call_expr)
	mut is_option := t.expr_returns_option(call_expr)

	// Fallback to function name lookup for simple function calls
	fn_name := t.get_call_fn_name(call_expr)
	if !is_result && !is_option && fn_name != '' {
		is_result = t.fn_returns_result(fn_name)
		is_option = t.fn_returns_option(fn_name)
	}

	if !is_result && !is_option {
		// V only allows `or` on Result/Option expressions.
		// If type lookup fails, default to Result (more common).
		is_result = true
	}

	// Native backends (arm64/x64) don't use Option/Result structs.
	// Expand `fn() or { fallback }` to: { _t := fn(); if _t { _t } else { fallback } }
	if t.pref != unsafe { nil } && (t.pref.backend == .arm64 || t.pref.backend == .x64) {
		temp_name := t.gen_temp_name()
		temp_ident := ast.Ident{
			name: temp_name
		}
		// For ?SumType returns, use _data field check instead of raw truthiness.
		mut base_type_name2 := t.get_expr_base_type(call_expr)
		if base_type_name2 == '' {
			if fn_name != '' {
				base_type_name2 = t.get_fn_return_base_type(fn_name)
			}
		}
		is_sumtype_return2 := base_type_name2 != '' && t.is_sum_type(base_type_name2)
		synth_pos3 := t.next_synth_pos()
		cond_expr2 := if is_sumtype_return2 {
			t.synth_selector(temp_ident, '_data', types.Type(types.voidptr_))
		} else {
			ast.Expr(temp_ident)
		}
		not_cond_expr2 := if is_sumtype_return2 {
			ast.Expr(ast.PrefixExpr{
				op:   .not
				expr: t.synth_selector(ast.Ident{
					name: temp_name
					pos:  synth_pos3
				}, '_data', types.Type(types.voidptr_))
			})
		} else {
			ast.Expr(ast.PrefixExpr{
				op:   .not
				expr: temp_ident
			})
		}
		prefix_stmts << ast.AssignStmt{
			op:  .decl_assign
			lhs: [ast.Expr(temp_ident)]
			rhs: [t.transform_expr(call_expr)]
		}
		or_side_effect_stmts, or_value := t.get_or_block_stmts_and_value(or_expr.stmts)
		// If there are side-effect statements, wrap in: if !_t._data { side_effects... }
		if or_side_effect_stmts.len > 0 {
			prefix_stmts << ast.ExprStmt{
				expr: ast.IfExpr{
					cond:  not_cond_expr2
					stmts: or_side_effect_stmts
				}
			}
		}
		return ast.IfExpr{
			cond:      cond_expr2
			stmts:     [ast.Stmt(ast.ExprStmt{
				expr: temp_ident
			})]
			else_expr: or_value
		}
	}

	// Get base type using expression-based lookup first, then fallback
	mut base_type := t.get_expr_base_type(call_expr)
	if base_type == '' && fn_name != '' {
		base_type = t.get_fn_return_base_type(fn_name)
	}
	// Generate temp variable name
	temp_name := t.gen_temp_name()
	temp_ident := ast.Ident{
		name: temp_name
	}
	if call_type := t.get_expr_type(call_expr) {
		if call_type is types.OptionType || call_type is types.ResultType {
			t.register_temp_var(temp_name, call_type)
			// Correct is_result/is_option based on resolved type
			if call_type is types.OptionType {
				is_result = false
				is_option = true
			} else if call_type is types.ResultType {
				is_result = true
				is_option = false
			}
			if base_type == '' {
				if call_type is types.ResultType {
					base_type = call_type.base_type.name()
				} else if call_type is types.OptionType {
					base_type = call_type.base_type.name()
				}
			}
		} else if ret_type := t.get_method_return_type(call_expr) {
			if ret_type is types.OptionType || ret_type is types.ResultType {
				t.register_temp_var(temp_name, ret_type)
				if ret_type is types.OptionType {
					is_result = false
					is_option = true
				} else if ret_type is types.ResultType {
					is_result = true
					is_option = false
				}
				if base_type == '' {
					if ret_type is types.ResultType {
						base_type = ret_type.base_type.name()
					} else if ret_type is types.OptionType {
						base_type = ret_type.base_type.name()
					}
				}
			}
		} else if fn_name != '' {
			if fn_ret := t.get_fn_return_type(fn_name) {
				if fn_ret is types.OptionType || fn_ret is types.ResultType {
					t.register_temp_var(temp_name, fn_ret)
					if fn_ret is types.OptionType {
						is_result = false
						is_option = true
					} else if fn_ret is types.ResultType {
						is_result = true
						is_option = false
					}
					if base_type == '' {
						if fn_ret is types.ResultType {
							base_type = fn_ret.base_type.name()
						} else if fn_ret is types.OptionType {
							base_type = fn_ret.base_type.name()
						}
					}
				}
			}
		}
	} else {
		if ret_type := t.get_method_return_type(call_expr) {
			// Fallback: get_expr_type may fail for method calls on complex expressions
			// (e.g. slices) where the checker didn't store a type at the call position.
			// Use get_method_return_type which resolves the receiver type and looks up
			// the method in the environment.
			t.register_temp_var(temp_name, ret_type)
			// Correct is_result/is_option based on resolved type
			if ret_type is types.OptionType {
				is_result = false
				is_option = true
			} else if ret_type is types.ResultType {
				is_result = true
				is_option = false
			}
			if base_type == '' {
				if ret_type is types.ResultType {
					base_type = ret_type.base_type.name()
				} else if ret_type is types.OptionType {
					base_type = ret_type.base_type.name()
				}
			}
		}
	}
	if base_type == '' && (is_result || is_option) {
		base_type = 'int'
	}
	// String range or-block: register as _result_string since the checker
	// didn't record a Result type for this expression.
	if is_string_range_or {
		t.register_temp_var(temp_name, types.ResultType{
			base_type: types.string_
		})
		base_type = 'string'
	}
	is_void_result := base_type == '' || base_type == 'void'
	// 1. _t1 := call_expr
	transformed_call2 := t.transform_expr(call_expr)
	// For string range or-blocks, rename string__substr to string__substr_with_check
	// which returns !string (Result) instead of string.
	rhs_expr2 := if is_string_range_or {
		t.rename_substr_to_checked(transformed_call2)
	} else {
		transformed_call2
	}
	prefix_stmts << ast.AssignStmt{
		op:  .decl_assign
		lhs: [ast.Expr(temp_ident)]
		rhs: [rhs_expr2]
	}
	// 2. if _t1.is_error { ... } (for Result) or if _t1.state != 0 { ... } (for Option)
	error_cond := if is_result {
		// _t1.is_error
		t.synth_selector(temp_ident, 'is_error', types.Type(types.bool_))
	} else {
		// _t1.state != 0
		ast.Expr(ast.InfixExpr{
			op:  .ne
			lhs: t.synth_selector(temp_ident, 'state', types.Type(types.int_))
			rhs: ast.BasicLiteral{
				kind:  .number
				value: '0'
			}
		})
	}
	// Build the if-block statements
	mut if_stmts := []ast.Stmt{}
	// Keep `err` available in or-block expansions; transformed interpolation
	// paths can reference it after this pass.
	if_stmts << ast.AssignStmt{
		op:  .decl_assign
		lhs: [ast.Expr(ast.Ident{
			name: 'err'
		})]
		rhs: [
			t.synth_selector(temp_ident, 'err', types.Type(types.Struct{
				name: 'IError'
			})),
		]
	}
	// Check if or-block contains a return statement (control flow)
	if t.or_block_has_return(or_expr.stmts) {
		// Or-block contains return - transform statements here to handle string
		// concatenation and other transformations. This is done here instead of
		// relying on later transform_stmt to avoid double smartcast transformation.
		if_stmts << t.transform_stmts(or_expr.stmts)
	} else if !is_void_result {
		// Or-block provides a value - assign to data (only for non-void results)
		or_side_effect_stmts, or_value := t.get_or_block_stmts_and_value(or_expr.stmts)
		if or_side_effect_stmts.len > 0 {
			if_stmts << or_side_effect_stmts
		}
		// Check if or-value is a void function call (e.g. error_with_pos()).
		// Void calls can't be assigned - treat as control flow instead.
		if t.is_void_call_expr(or_value) {
			if_stmts << ast.ExprStmt{
				expr: or_value
			}
		} else {
			// _t1.data = or_value
			if_stmts << ast.AssignStmt{
				op:  .assign
				lhs: [
					t.synth_selector(temp_ident, 'data', types.Type(types.voidptr_)),
				]
				rhs: [or_value]
			}
		}
	}
	prefix_stmts << ast.ExprStmt{
		expr: ast.IfExpr{
			cond:  error_cond
			stmts: if_stmts
		}
	}
	// Return the data access expression (or empty expr for void)
	if is_void_result {
		// For void results, return an empty expression since there's no value
		return ast.empty_expr
	}
	return t.synth_selector(temp_ident, 'data', types.Type(types.voidptr_))
}

// typed_deref generates a typed dereference of a voidptr:
// *unsafe { &ValueType(ptr) }
// This is needed because map__get_check returns voidptr, and dereferencing
// voidptr in the SSA builder loads only 1 byte (i8). The typed deref
// emits bitcast(ptr, *ValueType) + load(*ValueType) for correct load size.
fn (t &Transformer) typed_deref(ptr ast.Expr, value_type types.Type) ast.Expr {
	// For native backends (arm64/x64), map__get_check returns voidptr and
	// dereferencing voidptr loads only 1 byte (i8). Emit bitcast to correct
	// pointer type first: *(&ValueType(ptr))
	is_native := t.pref != unsafe { nil } && (t.pref.backend == .arm64 || t.pref.backend == .x64)
	if is_native {
		type_name := t.type_to_name(value_type)
		if type_name != '' {
			return ast.PrefixExpr{
				op:   .mul
				expr: ast.PrefixExpr{
					op:   .amp
					expr: ast.CastExpr{
						typ:  ast.Ident{
							name: type_name
						}
						expr: ptr
					}
				}
			}
		}
	}
	// C/cleanc backends handle voidptr deref correctly via C casts
	return ast.PrefixExpr{
		op:   .mul
		expr: ptr
	}
}

// try_expand_map_index_or handles the pattern: map[key] or { fallback }
// Transforms it to use map_get_check for safe lookup with fallback.
// Returns none if not a map index expression.
fn (mut t Transformer) try_expand_map_index_or(or_expr ast.OrExpr, mut prefix_stmts []ast.Stmt) ?ast.Expr {
	// Check if the inner expression is an IndexExpr
	if or_expr.expr !is ast.IndexExpr {
		return none
	}
	index_expr := or_expr.expr as ast.IndexExpr

	// Get the map type from environment and extract key/value types
	map_expr_typ := t.get_expr_type(index_expr.lhs) or { return none }
	map_type := t.unwrap_map_type(map_expr_typ) or { return none }
	value_type := map_type.value_type

	// Generate temp variable name for the pointer result
	temp_name := t.gen_temp_name()
	temp_ident := ast.Ident{
		name: temp_name
	}

	// Register temp variable type: get_check returns pointer to value type
	pointer_type := types.Pointer{
		base_type: value_type
	}
	t.register_temp_var(temp_name, pointer_type)

	map_arg := if t.is_pointer_type(map_expr_typ) {
		t.transform_expr(index_expr.lhs)
	} else {
		t.addr_of_expr_with_temp(index_expr.lhs, map_expr_typ)
	}

	// 1. Generate: _t1 := map__get_check(&m, &key)
	// This returns a pointer to the value, or null if not found
	get_check_call := ast.CallExpr{
		lhs:  ast.Ident{
			name: 'map__get_check'
		}
		args: [
			map_arg,
			t.voidptr_cast(t.addr_of_expr_with_temp(index_expr.expr, map_type.key_type)),
		]
	}
	prefix_stmts << ast.AssignStmt{
		op:  .decl_assign
		lhs: [ast.Expr(temp_ident)]
		rhs: [ast.Expr(get_check_call)]
	}

	// Check if or block has control flow (return/break/continue)
	has_control_flow := t.or_block_has_return(or_expr.stmts)

	// 2. Generate: if _t1 == nil { ... }
	null_check := ast.InfixExpr{
		op:  .eq
		lhs: temp_ident
		rhs: ast.Ident{
			name: 'nil'
		}
	}

	if has_control_flow {
		// Or block has control flow - use the statements directly
		// The control flow will exit, so we just dereference after
		prefix_stmts << ast.ExprStmt{
			expr: ast.IfExpr{
				cond:  null_check
				stmts: t.transform_stmts(or_expr.stmts)
			}
		}
	} else {
		// Or block provides a fallback value
		// We use two statements:
		// 1. result := fallback
		// 2. if ptr != nil { result = *ptr }
		result_temp := t.gen_temp_name()
		result_ident := ast.Ident{
			name: result_temp
		}

		// Register result temp variable with value type (not pointer)
		t.register_temp_var(result_temp, value_type)

		// Declare result with fallback value
		prefix_stmts << ast.AssignStmt{
			op:  .decl_assign
			lhs: [ast.Expr(result_ident)]
			rhs: [t.get_or_block_value(or_expr.stmts)]
		}

		// If ptr != nil, overwrite with actual value
		prefix_stmts << ast.ExprStmt{
			expr: ast.IfExpr{
				cond:  ast.InfixExpr{
					op:  .ne
					lhs: temp_ident
					rhs: ast.Ident{
						name: 'nil'
					}
				}
				stmts: [
					ast.Stmt(ast.AssignStmt{
						op:  .assign
						lhs: [ast.Expr(result_ident)]
						rhs: [t.typed_deref(temp_ident, value_type)]
					}),
				]
			}
		}
		return ast.Expr(result_ident)
	}

	// For control flow case, return the dereferenced pointer
	// (we know it's non-null because control flow would have exited)
	return t.typed_deref(temp_ident, value_type)
}

// try_expand_map_index_or_assign handles: var := map[key] or { fallback }
// Returns a list of statements that expand the assignment with proper map lookup.
fn (mut t Transformer) try_expand_map_index_or_assign(stmt ast.AssignStmt, or_expr ast.OrExpr) ?[]ast.Stmt {
	// Check if the inner expression is an IndexExpr
	if or_expr.expr !is ast.IndexExpr {
		return none
	}
	index_expr := or_expr.expr as ast.IndexExpr

	// Get the map type from environment and extract key/value types
	map_expr_typ := t.get_expr_type(index_expr.lhs) or { return none }
	map_type := t.unwrap_map_type(map_expr_typ) or { return none }
	value_type := map_type.value_type

	// Get the LHS variable name from the assignment
	if stmt.lhs.len != 1 {
		return none
	}

	mut stmts := []ast.Stmt{}

	// Generate temp variable name for the pointer result
	temp_name := t.gen_temp_name()
	temp_ident := ast.Ident{
		name: temp_name
	}

	// Register temp variable type: get_check returns pointer to value type
	pointer_type := types.Pointer{
		base_type: value_type
	}
	t.register_temp_var(temp_name, pointer_type)

	map_arg := if t.is_pointer_type(map_expr_typ) {
		t.transform_expr(index_expr.lhs)
	} else {
		t.addr_of_expr_with_temp(index_expr.lhs, map_expr_typ)
	}

	// 1. Generate: _t1 := map__get_check(&m, &key)
	get_check_call := ast.CallExpr{
		lhs:  ast.Ident{
			name: 'map__get_check'
		}
		args: [
			map_arg,
			t.voidptr_cast(t.addr_of_expr_with_temp(index_expr.expr, map_type.key_type)),
		]
	}
	stmts << ast.AssignStmt{
		op:  .decl_assign
		lhs: [ast.Expr(temp_ident)]
		rhs: [ast.Expr(get_check_call)]
		pos: stmt.pos
	}

	// Check if or block has control flow (return/break/continue)
	has_control_flow := t.or_block_has_return(or_expr.stmts)

	if has_control_flow {
		// Check if or block contains a nested map or block that needs expansion
		// e.g., scopes[k1] or { scopes[k2] or { return -999 } }
		mut has_nested_or := false
		for or_stmt in or_expr.stmts {
			if or_stmt is ast.ExprStmt {
				if or_stmt.expr is ast.OrExpr {
					inner_or := or_stmt.expr as ast.OrExpr
					if inner_or.expr is ast.IndexExpr {
						has_nested_or = true
						break
					}
				}
			}
		}

		if has_nested_or {
			// For nested or blocks, we need to declare the outer variable first
			// so we can assign to it inside the nested expansion
			// Pattern:
			// 1. lhs := 0 (default)
			// 2. if ptr1 == nil { ... nested ... lhs = nested_result }
			// 3. if ptr1 != nil { lhs = *ptr1 }

			// 1. Declare lhs with zero value
			stmts << ast.AssignStmt{
				op:  stmt.op
				lhs: stmt.lhs
				rhs: [
					ast.Expr(ast.BasicLiteral{
						kind:  .number
						value: '0'
					}),
				]
				pos: stmt.pos
			}

			// 2. Expand the nested or block in the null case
			null_check := ast.InfixExpr{
				op:  .eq
				lhs: temp_ident
				rhs: ast.Ident{
					name: 'nil'
				}
			}
			mut expanded_or_stmts := []ast.Stmt{}
			for or_stmt in or_expr.stmts {
				if or_stmt is ast.ExprStmt {
					expr_stmt := or_stmt as ast.ExprStmt
					if expr_stmt.expr is ast.OrExpr {
						inner_or := expr_stmt.expr as ast.OrExpr
						if inner_or.expr is ast.IndexExpr {
							// Create an assignment for the nested or
							inner_assign := ast.AssignStmt{
								op:  .assign
								lhs: stmt.lhs
								rhs: [ast.Expr(inner_or)]
							}
							if inner_stmts := t.try_expand_map_index_or_assign(inner_assign,
								inner_or)
							{
								expanded_or_stmts << inner_stmts
								continue
							}
						}
					}
				}
				expanded_or_stmts << or_stmt
			}
			stmts << ast.ExprStmt{
				expr: ast.IfExpr{
					cond:  null_check
					stmts: expanded_or_stmts
				}
			}

			// 3. If outer lookup succeeded, assign deref
			stmts << ast.ExprStmt{
				expr: ast.IfExpr{
					cond:  ast.InfixExpr{
						op:  .ne
						lhs: temp_ident
						rhs: ast.Ident{
							name: 'nil'
						}
					}
					stmts: [
						ast.Stmt(ast.AssignStmt{
							op:  .assign
							lhs: stmt.lhs
							rhs: [t.typed_deref(temp_ident, value_type)]
						}),
					]
				}
			}
		} else {
			// Simple control flow case (e.g., return inside or block)
			null_check := ast.InfixExpr{
				op:  .eq
				lhs: temp_ident
				rhs: ast.Ident{
					name: 'nil'
				}
			}
			stmts << ast.ExprStmt{
				expr: ast.IfExpr{
					cond:  null_check
					stmts: t.transform_stmts(or_expr.stmts)
				}
			}
			// lhs := *_t1 (typed deref for correct load size)
			stmts << ast.AssignStmt{
				op:  stmt.op
				lhs: stmt.lhs
				rhs: [t.typed_deref(temp_ident, value_type)]
				pos: stmt.pos
			}
		}
	} else {
		// 2b. lhs := fallback
		stmts << ast.AssignStmt{
			op:  stmt.op
			lhs: stmt.lhs
			rhs: [t.get_or_block_value(or_expr.stmts)]
			pos: stmt.pos
		}
		// 3b. if _t1 != nil { lhs = *_t1 } (typed deref for correct load size)
		stmts << ast.ExprStmt{
			expr: ast.IfExpr{
				cond:  ast.InfixExpr{
					op:  .ne
					lhs: temp_ident
					rhs: ast.Ident{
						name: 'nil'
					}
				}
				stmts: [
					ast.Stmt(ast.AssignStmt{
						op:  .assign
						lhs: stmt.lhs
						rhs: [t.typed_deref(temp_ident, value_type)]
					}),
				]
			}
		}
	}

	return stmts
}

// shared_mtx_expr creates the mutex access expression for a shared variable.
// For struct field access (e.g., e.scores), use the parent object's .mtx => e.mtx
// For standalone variables (e.g., data), use data.mtx
fn (mut t Transformer) shared_mtx_expr(locked_expr ast.Expr) ast.Expr {
	if locked_expr is ast.SelectorExpr {
		// Struct field: e.scores => e.mtx
		return t.synth_selector(locked_expr.lhs, 'mtx', types.Type(types.Struct{
			name: 'sync__RwMutex'
		}))
	}
	// Standalone variable: data => data.mtx
	return t.synth_selector(locked_expr, 'mtx', types.Type(types.Struct{
		name: 'sync__RwMutex'
	}))
}

// expand_lock_expr lowers a LockExpr into mutex lock/unlock calls around the body.
// lock data { body } => sync__RwMutex_lock(&data.mtx); body; sync__RwMutex_unlock(&data.mtx);
// rlock data { body } => sync__RwMutex_rlock(&data.mtx); body; sync__RwMutex_runlock(&data.mtx);
fn (mut t Transformer) expand_lock_expr(expr ast.LockExpr) []ast.Stmt {
	mut result := []ast.Stmt{}
	// For native backends (arm64/x64), skip lock/unlock calls since there's
	// no threading support and the sync module is not available.
	is_native := t.pref != unsafe { nil } && (t.pref.backend == .arm64 || t.pref.backend == .x64)
	// Emit lock calls
	if !is_native {
		for lock_expr in expr.lock_exprs {
			result << ast.ExprStmt{
				expr: ast.CallExpr{
					lhs:  ast.Ident{
						name: 'sync__RwMutex_lock'
					}
					args: [
						ast.Expr(ast.PrefixExpr{
							op:   .amp
							expr: t.shared_mtx_expr(lock_expr)
						}),
					]
				}
			}
		}
		// Emit rlock calls
		for rlock_expr in expr.rlock_exprs {
			result << ast.ExprStmt{
				expr: ast.CallExpr{
					lhs:  ast.Ident{
						name: 'sync__RwMutex_rlock'
					}
					args: [
						ast.Expr(ast.PrefixExpr{
							op:   .amp
							expr: t.shared_mtx_expr(rlock_expr)
						}),
					]
				}
			}
		}
	}
	// Emit transformed body stmts
	for stmt in t.transform_stmts(expr.stmts) {
		result << stmt
	}
	// Emit unlock calls (reverse order of lock)
	if !is_native {
		for lock_expr in expr.lock_exprs {
			result << ast.ExprStmt{
				expr: ast.CallExpr{
					lhs:  ast.Ident{
						name: 'sync__RwMutex_unlock'
					}
					args: [
						ast.Expr(ast.PrefixExpr{
							op:   .amp
							expr: t.shared_mtx_expr(lock_expr)
						}),
					]
				}
			}
		}
		// Emit runlock calls (reverse order of rlock)
		for rlock_expr in expr.rlock_exprs {
			result << ast.ExprStmt{
				expr: ast.CallExpr{
					lhs:  ast.Ident{
						name: 'sync__RwMutex_runlock'
					}
					args: [
						ast.Expr(ast.PrefixExpr{
							op:   .amp
							expr: t.shared_mtx_expr(rlock_expr)
						}),
					]
				}
			}
		}
	}
	return result
}

// lower_defer_stmts collects DeferStmts from the function body (at any nesting level),
// removes them, and injects their bodies before every return statement (and at the end
// of the function). Defers execute in LIFO order (last defer first).
fn (mut t Transformer) lower_defer_stmts(stmts []ast.Stmt, has_return_type bool) []ast.Stmt {
	if !t.has_defer_stmt(stmts) {
		return stmts
	}
	// Lower defers in source order so returns before a defer do not run it.
	mut active_defers := [][]ast.Stmt{}
	mut lowered := t.lower_defer_block(stmts, mut active_defers, has_return_type)
	if lowered.len == 0 || !t.stmt_ends_with_return(lowered[lowered.len - 1]) {
		t.append_defer_bodies(mut lowered, active_defers)
	}
	return lowered
}

fn (t &Transformer) has_defer_stmt(stmts []ast.Stmt) bool {
	for stmt in stmts {
		match stmt {
			ast.DeferStmt {
				return true
			}
			ast.ExprStmt {
				if stmt.expr is ast.IfExpr {
					if t.has_defer_stmt(stmt.expr.stmts) {
						return true
					}
					if stmt.expr.else_expr is ast.IfExpr {
						if t.has_defer_stmt(stmt.expr.else_expr.stmts) {
							return true
						}
					}
				} else if stmt.expr is ast.UnsafeExpr {
					if t.has_defer_stmt(stmt.expr.stmts) {
						return true
					}
				}
			}
			ast.ForStmt {
				if t.has_defer_stmt(stmt.stmts) {
					return true
				}
			}
			ast.BlockStmt {
				if t.has_defer_stmt(stmt.stmts) {
					return true
				}
			}
			else {}
		}
	}
	return false
}

fn (mut t Transformer) append_defer_bodies(mut out []ast.Stmt, defer_bodies [][]ast.Stmt) {
	for i := defer_bodies.len - 1; i >= 0; i-- {
		out << defer_bodies[i]
	}
}

fn (t &Transformer) copy_defer_stack(active_defers [][]ast.Stmt) [][]ast.Stmt {
	mut copied := [][]ast.Stmt{cap: active_defers.len}
	for defer_body in active_defers {
		mut body_copy := []ast.Stmt{cap: defer_body.len}
		for stmt in defer_body {
			body_copy << stmt
		}
		copied << body_copy
	}
	return copied
}

fn (mut t Transformer) lower_defer_else(else_expr ast.Expr, active_defers [][]ast.Stmt, has_return_type bool) ast.Expr {
	if else_expr is ast.IfExpr {
		mut branch_defers := t.copy_defer_stack(active_defers)
		return ast.IfExpr{
			cond:      else_expr.cond
			stmts:     t.lower_defer_block(else_expr.stmts, mut branch_defers, has_return_type)
			else_expr: t.lower_defer_else(else_expr.else_expr, active_defers, has_return_type)
		}
	}
	return else_expr
}

fn (mut t Transformer) lower_defer_block(stmts []ast.Stmt, mut active_defers [][]ast.Stmt, has_return_type bool) []ast.Stmt {
	mut result := []ast.Stmt{cap: stmts.len}
	for stmt in stmts {
		match stmt {
			ast.DeferStmt {
				active_defers << stmt.stmts
			}
			ast.ReturnStmt {
				if active_defers.len == 0 {
					result << ast.Stmt(stmt)
				} else if has_return_type && stmt.exprs.len > 0 {
					t.temp_counter++
					temp_name := '_defer_t${t.temp_counter}'
					if expr_type := t.get_expr_type(stmt.exprs[0]) {
						t.register_temp_var(temp_name, expr_type)
					}
					ret_expr := ast.Expr(stmt.exprs[0])
					result << ast.Stmt(ast.AssignStmt{
						op:  .decl_assign
						lhs: [ast.Expr(ast.Ident{
							name: temp_name
						})]
						rhs: [ret_expr]
					})
					t.append_defer_bodies(mut result, active_defers)
					result << ast.Stmt(ast.ReturnStmt{
						exprs: [ast.Expr(ast.Ident{
							name: temp_name
						})]
					})
				} else {
					t.append_defer_bodies(mut result, active_defers)
					result << ast.Stmt(stmt)
				}
			}
			ast.ExprStmt {
				if stmt.expr is ast.IfExpr {
					mut then_defers := t.copy_defer_stack(active_defers)
					result << ast.Stmt(ast.ExprStmt{
						expr: ast.IfExpr{
							cond:      stmt.expr.cond
							stmts:     t.lower_defer_block(stmt.expr.stmts, mut then_defers,
								has_return_type)
							else_expr: t.lower_defer_else(stmt.expr.else_expr, active_defers,
								has_return_type)
						}
					})
				} else if stmt.expr is ast.UnsafeExpr {
					mut unsafe_defers := t.copy_defer_stack(active_defers)
					result << ast.Stmt(ast.ExprStmt{
						expr: ast.UnsafeExpr{
							stmts: t.lower_defer_block(stmt.expr.stmts, mut unsafe_defers,
								has_return_type)
						}
					})
				} else {
					result << ast.Stmt(stmt)
				}
			}
			ast.ForStmt {
				mut loop_defers := t.copy_defer_stack(active_defers)
				result << ast.Stmt(ast.ForStmt{
					init:  stmt.init
					cond:  stmt.cond
					post:  stmt.post
					stmts: t.lower_defer_block(stmt.stmts, mut loop_defers, has_return_type)
				})
			}
			ast.BlockStmt {
				mut block_defers := t.copy_defer_stack(active_defers)
				result << ast.Stmt(ast.BlockStmt{
					stmts: t.lower_defer_block(stmt.stmts, mut block_defers, has_return_type)
				})
			}
			else {
				result << stmt
			}
		}
	}
	return result
}

// collect_and_remove_defers recursively walks statements, collects DeferStmt bodies,
// and returns the statements with DeferStmts removed.
fn (mut t Transformer) collect_and_remove_defers(stmts []ast.Stmt, mut defer_bodies [][]ast.Stmt) []ast.Stmt {
	mut result := []ast.Stmt{cap: stmts.len}
	for stmt in stmts {
		match stmt {
			ast.DeferStmt {
				defer_bodies << stmt.stmts
			}
			ast.ExprStmt {
				expr := stmt.expr
				if expr is ast.IfExpr {
					cleaned_if := t.collect_defers_in_if(expr, mut defer_bodies)
					result << ast.Stmt(ast.ExprStmt{
						expr: cleaned_if
					})
				} else if expr is ast.UnsafeExpr {
					cleaned_stmts := t.collect_and_remove_defers(expr.stmts, mut defer_bodies)
					result << ast.Stmt(ast.ExprStmt{
						expr: ast.UnsafeExpr{
							stmts: cleaned_stmts
						}
					})
				} else {
					result << ast.Stmt(stmt)
				}
			}
			ast.ForStmt {
				result << ast.Stmt(ast.ForStmt{
					init:  stmt.init
					cond:  stmt.cond
					post:  stmt.post
					stmts: t.collect_and_remove_defers(stmt.stmts, mut defer_bodies)
				})
			}
			ast.BlockStmt {
				result << ast.Stmt(ast.BlockStmt{
					stmts: t.collect_and_remove_defers(stmt.stmts, mut defer_bodies)
				})
			}
			else {
				result << stmt
			}
		}
	}
	return result
}

fn (t &Transformer) stmt_ends_with_return(stmt ast.Stmt) bool {
	return stmt is ast.ReturnStmt
}

fn (mut t Transformer) transform_return_stmt(stmt ast.ReturnStmt) ast.ReturnStmt {
	// Native backends (arm64/x64) don't use Option/Result structs.
	// `return error(...)` and `return none` should be lowered to `return 0` (error/none indicator).
	if t.pref != unsafe { nil } && (t.pref.backend == .arm64 || t.pref.backend == .x64) {
		error_fn_names := ['error', 'error_posix', 'error_with_code', 'error_win32']
		if stmt.exprs.len == 1 {
			ret_expr := stmt.exprs[0]
			// Check for `error(...)` / `error_posix(...)` call — appears as CallOrCastExpr with lhs=Ident
			if ret_expr is ast.CallOrCastExpr {
				if ret_expr.lhs is ast.Ident && ret_expr.lhs.name in error_fn_names {
					return ast.ReturnStmt{
						exprs: [
							ast.Expr(ast.BasicLiteral{
								kind:  .number
								value: '0'
							}),
						]
					}
				}
			}
			// Also check for CallExpr form
			if ret_expr is ast.CallExpr {
				if ret_expr.lhs is ast.Ident && ret_expr.lhs.name in error_fn_names {
					return ast.ReturnStmt{
						exprs: [
							ast.Expr(ast.BasicLiteral{
								kind:  .number
								value: '0'
							}),
						]
					}
				}
			}
			// Check for `return none` — appears as Ident{name:'none'}
			if ret_expr is ast.Ident && ret_expr.name == 'none' {
				return ast.ReturnStmt{
					exprs: [
						ast.Expr(ast.BasicLiteral{
							kind:  .number
							value: '0'
						}),
					]
				}
			}
		}
	}
	mut exprs := []ast.Expr{cap: stmt.exprs.len}
	for expr in stmt.exprs {
		// Resolve enum shorthands in return expressions (e.g., return .string → token__Token__string)
		if t.cur_fn_ret_type_name != '' {
			if expr is ast.SelectorExpr {
				sel := expr as ast.SelectorExpr
				if sel.lhs is ast.EmptyExpr {
					resolved := t.resolve_enum_shorthand(expr, t.cur_fn_ret_type_name)
					exprs << t.transform_expr(resolved)
					continue
				}
			}
		}
		// If the return expression is a MatchExpr and the return type is a sum type,
		// set sumtype_return_wrap so transform_match_expr wraps each branch value
		if expr is ast.MatchExpr && t.cur_fn_ret_type_name != ''
			&& t.is_sum_type(t.cur_fn_ret_type_name) {
			old_wrap := t.sumtype_return_wrap
			t.sumtype_return_wrap = t.cur_fn_ret_type_name
			transformed := t.transform_expr(expr)
			t.sumtype_return_wrap = old_wrap
			exprs << transformed
			continue
		}
		// Before transforming, check if the expression is a smartcasted identifier
		// that needs re-wrapping into the return sum type
		mut smartcast_variant := ''
		if t.cur_fn_ret_type_name != '' && t.is_sum_type(t.cur_fn_ret_type_name) {
			if expr is ast.Ident {
				if ctx := t.find_smartcast_for_expr(expr.name) {
					smartcast_variant = ctx.variant
				}
			}
		}
		transformed := t.transform_expr(expr)
		// Wrap variant values in sum type initialization if needed.
		// Use wrap_sumtype_value_transformed because the value is already transformed above.
		// Using wrap_sumtype_value would transform the value a second time, causing
		// double smartcast dereferences (e.g., ((T*)(((T*)(x._data._T))->_data._T))->field).
		if t.cur_fn_ret_type_name != '' && t.is_sum_type(t.cur_fn_ret_type_name) {
			if wrapped := t.wrap_sumtype_value_transformed(transformed, t.cur_fn_ret_type_name) {
				exprs << wrapped
				continue
			}
			// If wrapping failed but we have a smartcast context, use the variant from it
			if smartcast_variant != '' {
				if wrapped := t.build_sumtype_init(transformed, smartcast_variant, t.cur_fn_ret_type_name) {
					exprs << wrapped
					continue
				}
			}
		}
		exprs << transformed
	}
	return ast.ReturnStmt{
		exprs: exprs
	}
}

fn (t &Transformer) unwrap_assoc_expr(expr ast.Expr) ?ast.AssocExpr {
	match expr {
		ast.AssocExpr {
			return expr
		}
		ast.ParenExpr {
			return t.unwrap_assoc_expr(expr.expr)
		}
		ast.ModifierExpr {
			return t.unwrap_assoc_expr(expr.expr)
		}
		else {
			return none
		}
	}
}

fn (mut t Transformer) gen_assoc_temp_name() string {
	t.temp_counter++
	return '_assoc_t${t.temp_counter}'
}

fn (mut t Transformer) lower_assoc_expr(node ast.AssocExpr, take_addr bool) ast.Expr {
	// {base | field: val} -> unsafe { tmp := Type(base); tmp.field = val; tmp }
	// &{base | field: val} -> unsafe { tmp := Type(base); tmp.field = val; &tmp }
	mut target_c := ''
	if target_type := t.get_expr_type(ast.Expr(node)) {
		target_c = t.type_to_c_name(target_type)
	}
	tmp_name := t.gen_assoc_temp_name()
	tmp_ident := ast.Ident{
		name: tmp_name
		pos:  node.pos
	}

	// Prepare the base value for the update.
	mut base_value := t.transform_expr(node.expr)
	if base_type := t.get_expr_type(node.expr) {
		if base_type is types.SumType && target_c != '' {
			// Unwrap sum type variant for struct update: *((${T}*)sum._data._Tshort)
			ctx := SmartcastContext{
				expr:         ''
				variant:      target_c
				variant_full: target_c
				sumtype:      ''
			}
			base_value = t.apply_smartcast_direct_ctx(node.expr, ctx)
		} else if t.is_pointer_type(base_type) {
			base_value = ast.Expr(ast.PrefixExpr{
				op:   token.Token.mul
				expr: base_value
			})
		}
	}

	// Hoist temp declaration and field updates before current statement via pending_stmts.
	t.pending_stmts << ast.Stmt(ast.AssignStmt{
		op:  .decl_assign
		lhs: [ast.Expr(tmp_ident)]
		rhs: [
			ast.Expr(ast.CastExpr{
				typ:  node.typ
				expr: base_value
			}),
		]
		pos: node.pos
	})

	// Apply field updates.
	for field in node.fields {
		t.pending_stmts << ast.Stmt(ast.AssignStmt{
			op:  .assign
			lhs: [
				t.synth_selector_from_struct(tmp_ident, field.name, target_c),
			]
			rhs: [t.transform_expr(field.value)]
			pos: node.pos
		})
	}

	// Yield value or address.
	if take_addr {
		return ast.Expr(ast.PrefixExpr{
			op:   token.Token.amp
			expr: tmp_ident
		})
	}
	return ast.Expr(tmp_ident)
}

fn (t &Transformer) is_nil_expr(expr ast.Expr) bool {
	return match expr {
		ast.Ident {
			expr.name == 'nil'
		}
		ast.Keyword {
			expr.tok == .key_nil
		}
		ast.Type {
			expr is ast.NilType
		}
		ast.ParenExpr {
			t.is_nil_expr(expr.expr)
		}
		else {
			false
		}
	}
}

fn (t &Transformer) is_unsafe_nil_expr(expr ast.UnsafeExpr) bool {
	if expr.stmts.len != 1 {
		return false
	}
	stmt := expr.stmts[0]
	if stmt is ast.ExprStmt {
		return t.is_nil_expr(stmt.expr)
	}
	return false
}

fn (t &Transformer) can_take_address_expr(expr ast.Expr) bool {
	return match expr {
		ast.Ident, ast.SelectorExpr, ast.IndexExpr {
			true
		}
		// String literals compile to compound literals in C, which are addressable.
		// Using &(string){...} is safe and avoids statement-expression temporaries
		// whose address would escape scope when used as function call arguments.
		ast.StringLiteral, ast.InitExpr, ast.ArrayInitExpr {
			true
		}
		ast.PrefixExpr {
			expr.op == .mul
		}
		ast.ParenExpr {
			t.can_take_address_expr(expr.expr)
		}
		else {
			false
		}
	}
}

// addr_of_with_prefix_temp creates a &expr for addressable expressions, or emits a temp
// variable declaration into prefix_stmts and returns &tmp for non-addressable expressions.
// This avoids the scope-escape issue with UnsafeExpr temporaries in function call arguments.
fn (mut t Transformer) addr_of_with_prefix_temp(expr ast.Expr, typ types.Type, mut prefix_stmts []ast.Stmt) ast.Expr {
	transformed := t.transform_expr(expr)
	if t.can_take_address_expr(transformed) {
		return ast.PrefixExpr{
			op:   .amp
			expr: transformed
		}
	}
	tmp_name := t.gen_temp_name()
	tmp_ident := ast.Ident{
		name: tmp_name
	}
	t.register_temp_var(tmp_name, typ)
	prefix_stmts << ast.Stmt(ast.AssignStmt{
		op:  .decl_assign
		lhs: [ast.Expr(tmp_ident)]
		rhs: [transformed]
	})
	return ast.PrefixExpr{
		op:   .amp
		expr: ast.Expr(tmp_ident)
	}
}

fn (mut t Transformer) addr_of_expr_with_temp(expr ast.Expr, typ types.Type) ast.Expr {
	transformed := t.transform_expr(expr)
	if t.can_take_address_expr(transformed) {
		return ast.PrefixExpr{
			op:   .amp
			expr: transformed
		}
	}
	tmp_name := t.gen_temp_name()
	tmp_ident := ast.Ident{
		name: tmp_name
	}
	t.register_temp_var(tmp_name, typ)
	return ast.UnsafeExpr{
		stmts: [
			ast.Stmt(ast.AssignStmt{
				op:  .decl_assign
				lhs: [ast.Expr(tmp_ident)]
				rhs: [transformed]
			}),
			ast.Stmt(ast.ExprStmt{
				expr: ast.PrefixExpr{
					op:   .amp
					expr: ast.Expr(tmp_ident)
				}
			}),
		]
	}
}

fn (t &Transformer) voidptr_cast(expr ast.Expr) ast.Expr {
	return ast.Expr(ast.CastExpr{
		typ:  ast.Ident{
			name: 'voidptr'
		}
		expr: expr
	})
}

fn (mut t Transformer) lower_wrapper_payload_access(wrapper_expr ast.Expr, base_type_name string) ast.Expr {
	err_selector := t.synth_selector(wrapper_expr, 'err', types.Type(types.Struct{
		name: 'IError'
	}))
	addr_err := ast.PrefixExpr{
		op:   .amp
		expr: err_selector
	}
	u8_ptr := ast.CastExpr{
		typ:  ast.Ident{
			name: 'u8*'
		}
		expr: addr_err
	}
	payload_ptr := ast.InfixExpr{
		op:  .plus
		lhs: u8_ptr
		rhs: ast.KeywordOperator{
			op:    .key_sizeof
			exprs: [
				ast.Expr(ast.Ident{
					name: 'IError'
				}),
			]
		}
	}
	typed_ptr := ast.CastExpr{
		typ:  ast.Ident{
			name: '${base_type_name}*'
		}
		expr: payload_ptr
	}
	return ast.ParenExpr{
		expr: ast.PrefixExpr{
			op:   .mul
			expr: typed_ptr
		}
	}
}

fn (t &Transformer) get_sprintf_format_for_type(typ types.Type) string {
	match typ {
		types.String {
			return '%s'
		}
		types.Primitive {
			if typ.props.has(types.Properties.boolean) {
				return '%s'
			}
			if typ.props.has(types.Properties.float) {
				return '%f'
			}
			if typ.props.has(types.Properties.unsigned) {
				if typ.size == 64 {
					return '%llu'
				}
				return '%u'
			}
			// signed integers
			if typ.size == 64 {
				return '%lld'
			}
			return '%d'
		}
		types.Rune {
			return '%c'
		}
		types.Char {
			return '%c'
		}
		types.Enum {
			// Enums use their .str() method, so format is %s
			if _ := t.get_str_fn_name_for_type(typ) {
				return '%s'
			}
			return '%d'
		}
		types.Pointer {
			return '%p'
		}
		types.Alias {
			// For aliases to primitive types (e.g., ValueID = int),
			// use the base type's format directly.
			return t.get_sprintf_format_for_type(typ.base_type)
		}
		else {
			// Custom types (struct, array, map, sumtype) that have .str() methods
			if _ := t.get_str_fn_name_for_type(typ) {
				return '%s'
			}
			return '%d'
		}
	}
}

fn (mut t Transformer) resolve_sprintf_format(inter ast.StringInter) string {
	mut fmt := '%'
	if inter.width > 0 {
		fmt += '${inter.width}'
	}
	if inter.precision > 0 {
		fmt += '.${inter.precision}'
	}
	if inter.format != .unformatted {
		match inter.format {
			.decimal { fmt += 'd' }
			.float { fmt += 'f' }
			.hex { fmt += 'x' }
			.octal { fmt += 'o' }
			.character { fmt += 'c' }
			.exponent { fmt += 'e' }
			.exponent_short { fmt += 'g' }
			.binary { fmt += 'd' } // binary not supported in printf, fallback to decimal
			.pointer_address { fmt += 'p' }
			.string { fmt += 's' }
			.unformatted { fmt += 'd' }
		}
		return fmt
	}
	// Infer from expression type
	if typ := t.get_expr_type(inter.expr) {
		return t.get_sprintf_format_for_type(typ)
	}
	return '%d' // fallback
}

fn (mut t Transformer) transform_sprintf_arg(inter ast.StringInter) ast.Expr {
	transformed := t.transform_expr(inter.expr)
	typ := t.get_expr_type(inter.expr) or {
		return transformed // can't resolve type, pass as-is
	}
	// When an explicit format is specified, pass the expression as-is.
	// The user has explicitly chosen the format, so no wrapping is needed
	// (e.g., ${ptr:p} should pass the pointer directly, not call .str()).
	if inter.format != .unformatted {
		if inter.format == .string {
			// Explicit :s still needs .str access for V strings
			if typ is types.String {
				return t.synth_selector(transformed, 'str', types.Type(types.voidptr_))
			}
		}
		return transformed
	}
	match typ {
		types.String {
			// string -> expr.str (access C char* pointer for sprintf %s)
			return t.synth_selector(transformed, 'str', types.Type(types.voidptr_))
		}
		types.Primitive {
			if typ.props.has(types.Properties.boolean) {
				// bool -> if expr { "true" } else { "false" } (ternary for %s)
				return ast.Expr(ast.IfExpr{
					cond:      transformed
					stmts:     [
						ast.Stmt(ast.ExprStmt{
							expr: ast.Expr(ast.StringLiteral{
								kind:  .c
								value: '"true"'
							})
						}),
					]
					else_expr: ast.Expr(ast.StringLiteral{
						kind:  .c
						value: '"false"'
					})
					pos:       inter.expr.pos()
				})
			}
			// numeric primitives: pass as-is
			return transformed
		}
		types.Rune, types.Char {
			return transformed
		}
		types.Enum {
			// Enums should call their .str() method for string representation
			if str_fn_name := t.get_str_fn_name_for_type(typ) {
				str_call := ast.Expr(ast.CallExpr{
					lhs:  ast.Ident{
						name: str_fn_name
					}
					args: [transformed]
					pos:  inter.expr.pos()
				})
				return t.synth_selector(str_call, 'str', types.Type(types.voidptr_))
			}
			return transformed
		}
		types.Alias {
			// For aliases to primitives (e.g., ValueID = int),
			// handle based on the base type to avoid calling non-existent str() functions.
			base := typ.base_type
			match base {
				types.String {
					return t.synth_selector(transformed, 'str', types.Type(types.voidptr_))
				}
				types.Primitive {
					if base.props.has(types.Properties.boolean) {
						return ast.Expr(ast.IfExpr{
							cond:      transformed
							stmts:     [
								ast.Stmt(ast.ExprStmt{
									expr: ast.Expr(ast.StringLiteral{
										kind:  .c
										value: '"true"'
									})
								}),
							]
							else_expr: ast.Expr(ast.StringLiteral{
								kind:  .c
								value: '"false"'
							})
							pos:       inter.expr.pos()
						})
					}
					return transformed
				}
				else {
					return transformed
				}
			}
		}
		else {
			// For custom types with str() method: Type__str(expr).str
			str_fn_info := t.get_str_fn_info_for_expr(inter.expr)
			if str_fn_info.str_fn_name != '' {
				t.needed_str_fns[str_fn_info.str_fn_name] = str_fn_info.elem_type
				str_call := ast.Expr(ast.CallExpr{
					lhs:  ast.Ident{
						name: str_fn_info.str_fn_name
					}
					args: [transformed]
					pos:  inter.expr.pos()
				})
				return t.synth_selector(str_call, 'str', types.Type(types.voidptr_))
			}
			return transformed
		}
	}
}

fn (mut t Transformer) transform_string_inter_literal(expr ast.StringInterLiteral) ast.Expr {
	mut new_inters := []ast.StringInter{cap: expr.inters.len}
	for inter in expr.inters {
		new_inters << ast.StringInter{
			format:       inter.format
			width:        inter.width
			precision:    inter.precision
			expr:         t.transform_sprintf_arg(inter)
			format_expr:  inter.format_expr
			resolved_fmt: t.resolve_sprintf_format(inter)
		}
	}
	return ast.StringInterLiteral{
		kind:   expr.kind
		values: expr.values
		inters: new_inters
	}
}

// apply_smartcast_direct_ctx generates a cast expression for direct access to a smartcast variable
// For primitives: ((int)(intptr_t)v._data._int) - cast from pointer space back to value
// For structs/strings: (*((ast__Type*)v._data._Type)) - dereference pointer
fn (mut t Transformer) apply_smartcast_direct_ctx(original_expr ast.Expr, ctx SmartcastContext) ast.Expr {
	// variant (short name) is used for union member access: _data._Array_Attribute
	// variant_full (full name) is used for type cast: (Array_ast__Attribute*)
	variant_short := ctx.variant
	// Extract simple variant name for _data._ accessor (strip module prefix for non-composite types)
	// But preserve composite type prefixes like Array_, Map_, Array_fixed_
	variant_simple := if variant_short.starts_with('Array_') || variant_short.starts_with('Map_') {
		// For composite types (arrays, maps), use the short name to match union member
		variant_short
	} else if variant_short.contains('__') {
		variant_short.all_after_last('__')
	} else {
		variant_short
	}
	// For type cast, use the full variant name from context
	// This has the proper module prefix for the typedef
	mangled_variant := if ctx.variant_full != '' {
		ctx.variant_full
	} else if variant_short.contains('__') {
		variant_short // Already has module prefix
	} else if t.cur_module != '' && t.cur_module != 'main' && t.cur_module != 'builtin' {
		'${t.cur_module}__${variant_short}'
	} else {
		variant_short
	}
	// For nested smartcasts, transform the base expression first.
	// Temporarily remove this exact context to avoid applying it recursively.
	removed_ctxs := t.remove_matching_smartcasts(ctx)
	transformed_base := t.transform_expr(original_expr)
	t.restore_smartcasts(removed_ctxs)
	if t.expr_is_casted_to_type(transformed_base, '${mangled_variant}*') {
		return ast.ParenExpr{
			expr: ast.PrefixExpr{
				op:   token.Token.mul
				expr: transformed_base
			}
		}
	}
	// Already concretely casted to this variant by an outer smartcast context.
	if t.expr_is_casted_to_type(transformed_base, mangled_variant) {
		return transformed_base
	}
	// Create data access.
	// For native backends (arm64/x64): _data is a plain i64 (void pointer) in the SSA struct.
	// No union variant sub-field exists, so just use _data directly.
	// For C backends: _data is a union, so access _data._variant for the specific member.
	is_native_backend := t.pref != unsafe { nil }
		&& (t.pref.backend == .arm64 || t.pref.backend == .x64)
	data_access := t.synth_selector(transformed_base, '_data', types.Type(types.voidptr_))
	variant_access := if is_native_backend {
		data_access
	} else {
		t.synth_selector(data_access, '_${variant_simple}', types.Type(types.voidptr_))
	}

	// For primitives, cast from pointer space back to value type
	if variant_simple in ['int', 'i8', 'i16', 'i32', 'i64', 'u8', 'u16', 'u32', 'u64', 'f32', 'f64',
		'bool', 'rune', 'byte', 'usize', 'isize'] {
		// Create: ((variant)(intptr_t)variant_access)
		return ast.ParenExpr{
			expr: ast.CastExpr{
				typ:  ast.Ident{
					name: variant_simple
				}
				expr: ast.CastExpr{
					typ:  ast.Ident{
						name: 'intptr_t'
					}
					expr: variant_access
				}
			}
		}
	}

	// For structs/strings, dereference the pointer
	// Create: (mangled_variant*)variant_access
	cast_expr := ast.CastExpr{
		typ:  ast.Ident{
			name: '${mangled_variant}*'
		}
		expr: variant_access
	}
	// Create: *(cast_expr) wrapped in parens for proper precedence when accessing fields
	deref_expr := ast.PrefixExpr{
		op:   token.Token.mul
		expr: cast_expr
	}
	return ast.ParenExpr{
		expr: deref_expr
	}
}

// apply_smartcast_receiver_ctx generates a cast expression for a method call receiver on a smartcast variable
// e.g., se.lhs when smartcast to SelectorExpr -> (*((ast__SelectorExpr*)se.lhs._data._SelectorExpr))
fn (mut t Transformer) apply_smartcast_receiver_ctx(sumtype_expr ast.Expr, ctx SmartcastContext) ast.Expr {
	// variant (short name) is used for union member access
	// variant_full (full name) is used for type cast
	variant_short := ctx.variant
	// Extract simple variant name for _data._ accessor (strip module prefix)
	// But preserve composite type prefixes like Array_, Map_, Array_fixed_
	variant_simple := if variant_short.starts_with('Array_') || variant_short.starts_with('Map_') {
		// For composite types, use the short name to match union member
		variant_short
	} else if variant_short.contains('__') {
		variant_short.all_after_last('__')
	} else {
		variant_short
	}
	// Use full variant name for type cast from context
	mangled_variant := if ctx.variant_full != '' {
		ctx.variant_full
	} else if variant_short.contains('__') {
		variant_short // Already has module prefix
	} else if t.cur_module != '' && t.cur_module != 'main' && t.cur_module != 'builtin' {
		'${t.cur_module}__${variant_short}'
	} else {
		variant_short
	}
	// For nested smartcasts, transform the base expression first.
	// Temporarily remove this exact context to avoid applying it recursively.
	removed_ctxs := t.remove_matching_smartcasts(ctx)
	transformed_base := t.transform_expr(sumtype_expr)
	t.restore_smartcasts(removed_ctxs)
	if t.expr_is_casted_to_type(transformed_base, '${mangled_variant}*') {
		return ast.ParenExpr{
			expr: ast.PrefixExpr{
				op:   token.Token.mul
				expr: transformed_base
			}
		}
	}
	// Already concretely casted to this variant by an outer smartcast context.
	if t.expr_is_casted_to_type(transformed_base, mangled_variant) {
		return transformed_base
	}
	// Create data access.
	// For native backends: _data is a plain i64, no union variant sub-field.
	// For C backends: _data is a union, access _data._variant.
	is_native_backend2 := t.pref != unsafe { nil }
		&& (t.pref.backend == .arm64 || t.pref.backend == .x64)
	data_access := t.synth_selector(transformed_base, '_data', types.Type(types.voidptr_))
	variant_access := if is_native_backend2 {
		data_access
	} else {
		t.synth_selector(data_access, '_${variant_simple}', types.Type(types.voidptr_))
	}
	// Create: (mangled_variant*)variant_access
	cast_expr := ast.CastExpr{
		typ:  ast.Ident{
			name: '${mangled_variant}*'
		}
		expr: variant_access
	}
	// Create: *(cast_expr) - dereference to get the actual value
	deref_expr := ast.PrefixExpr{
		op:   token.Token.mul
		expr: cast_expr
	}
	return ast.ParenExpr{
		expr: deref_expr
	}
}

// apply_smartcast_field_access_ctx generates a cast expression for field access on a smartcast variable
// e.g., w.valera.name when smartcast to Kek -> ((ast__Kek*)w.valera._data._Kek)->name
// For nested smartcasts, we first transform the base expression to apply outer smartcasts

fn (mut t Transformer) build_match_branch_cond(match_expr ast.Expr, conds []ast.Expr, is_match_true bool, is_match_false bool) ast.Expr {
	mut branch_cond := ast.Expr(ast.empty_expr)
	for cond in conds {
		single_cond := t.build_single_match_cond(match_expr, cond, is_match_true, is_match_false)
		if branch_cond is ast.EmptyExpr {
			branch_cond = single_cond
		} else {
			branch_cond = ast.Expr(ast.InfixExpr{
				op:  .logical_or
				lhs: branch_cond
				rhs: single_cond
				pos: cond.pos()
			})
		}
	}
	return branch_cond
}

fn (mut t Transformer) build_single_match_cond(match_expr ast.Expr, cond ast.Expr, is_match_true bool, is_match_false bool) ast.Expr {
	if is_match_true || is_match_false {
		cond_expr := t.transform_expr(cond)
		if is_match_false {
			return ast.PrefixExpr{
				op:   .not
				expr: cond_expr
				pos:  cond.pos()
			}
		}
		return cond_expr
	}

	if cond is ast.RangeExpr {
		lower_bound := ast.InfixExpr{
			op:  .ge
			lhs: match_expr
			rhs: t.transform_expr(cond.start)
			pos: cond.pos
		}
		if cond.end is ast.EmptyExpr {
			return lower_bound
		}
		upper_op := if cond.op == .dotdot { token.Token.lt } else { token.Token.le }
		upper_bound := ast.InfixExpr{
			op:  upper_op
			lhs: match_expr
			rhs: t.transform_expr(cond.end)
			pos: cond.pos
		}
		return ast.InfixExpr{
			op:  .and
			lhs: lower_bound
			rhs: upper_bound
			pos: cond.pos
		}
	}

	return ast.InfixExpr{
		op:  .eq
		lhs: match_expr
		rhs: t.transform_expr(cond)
		pos: cond.pos()
	}
}

fn (t &Transformer) is_supported_struct_default_expr(expr ast.Expr) bool {
	match expr {
		ast.BasicLiteral, ast.StringLiteral, ast.SelectorExpr, ast.CallExpr, ast.CallOrCastExpr,
		ast.PrefixExpr, ast.CastExpr, ast.ArrayInitExpr, ast.MapInitExpr, ast.InitExpr {
			return true
		}
		ast.Ident {
			return expr.name !in ['none', 'none__']
		}
		else {
			return false
		}
	}
}

fn (t &Transformer) flatten_and_terms(expr ast.Expr) []ast.Expr {
	if expr is ast.InfixExpr && expr.op == token.Token.and {
		mut terms := []ast.Expr{}
		terms << t.flatten_and_terms(expr.lhs)
		terms << t.flatten_and_terms(expr.rhs)
		return terms
	}
	return [expr]
}

fn (t &Transformer) join_and_terms(terms []ast.Expr) ast.Expr {
	if terms.len == 0 {
		return ast.BasicLiteral{
			kind:  token.Token.key_true
			value: 'true'
		}
	}
	mut out := terms[0]
	for i in 1 .. terms.len {
		out = ast.Expr(ast.InfixExpr{
			op:  token.Token.and
			lhs: out
			rhs: terms[i]
		})
	}
	return out
}

fn (t &Transformer) smartcast_context_from_is_check(expr ast.InfixExpr) ?SmartcastContext {
	// checker can lower `is` into `.eq` with type RHS in some contexts.
	if expr.op !in [.key_is, .eq] {
		return none
	}
	mut variant_name := ''
	mut variant_module := ''
	if expr.rhs is ast.Ident {
		variant_name = (expr.rhs as ast.Ident).name
	} else if expr.rhs is ast.SelectorExpr {
		sel := expr.rhs as ast.SelectorExpr
		variant_name = sel.rhs.name
		if sel.lhs is ast.Ident {
			variant_module = (sel.lhs as ast.Ident).name
		}
	}
	if variant_name == '' {
		return none
	}
	if expr.op == .eq {
		lookup_name := if variant_module != '' {
			'${variant_module}__${variant_name}'
		} else {
			variant_name
		}
		if t.lookup_type(lookup_name) == none && t.lookup_type(variant_name) == none {
			return none
		}
	}

	mut sumtype_name := t.get_sumtype_name_for_expr(expr.lhs)
	if sumtype_name == '' {
		sumtype_name = t.find_sumtype_for_variant(variant_name)
	}
	if sumtype_name == '' {
		return none
	}

	variants := t.get_sum_type_variants(sumtype_name)
	mut has_variant := false
	mangled_variant := if variant_module != '' {
		'${variant_module}__${variant_name}'
	} else {
		variant_name
	}
	for v in variants {
		v_short := if v.contains('__') { v.all_after_last('__') } else { v }
		if v == variant_name || v_short == variant_name || v == mangled_variant
			|| v_short == mangled_variant {
			has_variant = true
			break
		}
	}
	if !has_variant {
		return none
	}

	qualified_variant := if variant_module != '' {
		'${variant_module}__${variant_name}'
	} else {
		variant_name
	}
	qualified_variant_full := if variant_module != '' {
		'${variant_module}__${variant_name}'
	} else if t.cur_module != '' && t.cur_module != 'main' && t.cur_module != 'builtin' {
		'${t.cur_module}__${variant_name}'
	} else {
		variant_name
	}
	return SmartcastContext{
		expr:         t.expr_to_string(expr.lhs)
		variant:      qualified_variant
		variant_full: qualified_variant_full
		sumtype:      sumtype_name
	}
}

// expr_to_string converts an expression to its string representation for smart cast matching
fn (t &Transformer) expr_to_string(expr ast.Expr) string {
	if expr is ast.Ident {
		return expr.name
	}
	if expr is ast.SelectorExpr {
		lhs_str := t.expr_to_string(expr.lhs)
		return '${lhs_str}.${expr.rhs.name}'
	}
	if expr is ast.ParenExpr {
		return t.expr_to_string(expr.expr)
	}
	if expr is ast.ModifierExpr {
		return t.expr_to_string(expr.expr)
	}
	return ''
}

// match_variant finds the variant in variants that matches c_name (exact or short name match)
fn (t &Transformer) match_variant(c_name string, variants []string) ?string {
	if c_name in variants {
		return c_name
	}
	c_short := if c_name.contains('__') { c_name.all_after_last('__') } else { c_name }
	for v in variants {
		v_short := if v.contains('__') { v.all_after_last('__') } else { v }
		if c_short == v_short || c_short == v {
			return v
		}
	}
	return none
}

fn (t &Transformer) is_array_value_expr(expr ast.Expr) bool {
	if t.get_array_elem_type_str(expr) != none {
		return true
	}
	if expr is ast.ParenExpr {
		return t.is_array_value_expr(expr.expr)
	}
	if expr is ast.PrefixExpr && expr.op == .mul {
		if t.get_array_elem_type_str(expr.expr) != none {
			return true
		}
		if inner_typ := t.get_expr_type(expr.expr) {
			if inner_typ is types.Pointer {
				mut base_typ := inner_typ.base_type
				if base_typ is types.Alias {
					base_typ = (base_typ as types.Alias).base_type
				}
				if base_typ is types.Array || base_typ is types.ArrayFixed {
					return true
				}
			}
		}
	}
	if typ := t.get_expr_type(expr) {
		mut base_typ := typ.base_type()
		if base_typ is types.Alias {
			base_typ = (base_typ as types.Alias).base_type
		}
		if base_typ is types.Array || base_typ is types.ArrayFixed {
			return true
		}
	}
	return false
}

fn (t &Transformer) get_array_method_info(expr ast.Expr) ?ArrayMethodInfo {
	if expr_type := t.get_expr_type(expr) {
		base_type := t.unwrap_alias_and_pointer_type(expr_type)
		match base_type {
			types.Array {
				elem_type_name := t.array_elem_type_name_for_helpers(base_type.elem_type)
				if elem_type_name == '' || elem_type_name == 'void' {
					return none
				}
				return ArrayMethodInfo{
					array_type: 'Array_${elem_type_name}'
					elem_type:  elem_type_name
					is_fixed:   false
				}
			}
			types.ArrayFixed {
				elem_type_name := t.array_elem_type_name_for_helpers(base_type.elem_type)
				if elem_type_name == '' || elem_type_name == 'void' {
					return none
				}
				return ArrayMethodInfo{
					array_type: 'Array_fixed_${elem_type_name}_${base_type.len}'
					elem_type:  elem_type_name
					is_fixed:   true
					fixed_len:  base_type.len
				}
			}
			else {}
		}
	}
	if arr_type := t.get_array_type_str(expr) {
		if arr_type.starts_with('Array_fixed_') {
			payload := arr_type['Array_fixed_'.len..]
			if payload.contains('_') {
				elem_type_name := payload.all_before_last('_')
				len_str := payload.all_after_last('_')
				if elem_type_name == '' || elem_type_name == 'void' {
					return none
				}
				return ArrayMethodInfo{
					array_type: arr_type
					elem_type:  elem_type_name
					is_fixed:   true
					fixed_len:  len_str.int()
				}
			}
		}
		if arr_type.starts_with('Array_') {
			elem_type_name := arr_type['Array_'.len..]
			if elem_type_name == '' || elem_type_name == 'void' {
				return none
			}
			return ArrayMethodInfo{
				array_type: arr_type
				elem_type:  elem_type_name
				is_fixed:   false
			}
		}
	}
	if elem_type_name := t.get_array_elem_type_str(expr) {
		if elem_type_name == '' || elem_type_name == 'void' {
			return none
		}
		return ArrayMethodInfo{
			array_type: 'Array_${elem_type_name}'
			elem_type:  elem_type_name
			is_fixed:   false
		}
	}
	return none
}

fn (mut t Transformer) register_needed_array_method(info ArrayMethodInfo, method_name string) string {
	fn_name := '${info.array_type}_${method_name}'
	match method_name {
		'contains' {
			t.needed_array_contains_fns[fn_name] = info
		}
		'index' {
			t.needed_array_index_fns[fn_name] = info
		}
		'last_index' {
			t.needed_array_last_index_fns[fn_name] = info
		}
		else {}
	}
	return fn_name
}

fn (mut t Transformer) transform_array_receiver_expr(receiver ast.Expr) ast.Expr {
	transformed := t.transform_expr(receiver)
	if recv_type := t.get_expr_type(receiver) {
		base_type := t.unwrap_alias_and_pointer_type(recv_type)
		if recv_type is types.Pointer && (base_type is types.Array || base_type is types.ArrayFixed) {
			return ast.PrefixExpr{
				op:   .mul
				expr: transformed
			}
		}
	}
	return transformed
}

// is_map_lookup_returning_array checks if an expression is a map lookup that returns an array type
fn (t &Transformer) is_map_lookup_returning_array(expr ast.Expr) bool {
	// Check if expr is an IndexExpr (map[key])
	if expr !is ast.IndexExpr {
		return false
	}
	index_expr := expr as ast.IndexExpr
	// Check if the LHS is a map type
	map_type := t.get_expr_type(index_expr.lhs) or { return false }
	if map_type is types.Map {
		// Check if the value type is an array
		return map_type.value_type is types.Array
	}
	return false
}

// transform_flag_enum_method transforms:
//   receiver.has(flag) → (int(receiver) & int(flag)) != 0
//   receiver.all(flags) → (int(receiver) & int(flags)) == int(flags)
fn (mut t Transformer) transform_flag_enum_method(receiver ast.Expr, method string, args []ast.Expr, enum_type string) ast.Expr {
	if args.len == 0 {
		return ast.empty_expr
	}

	arg := args[0]

	// Resolve enum shorthand: .read → EnumType__read
	resolved_arg := t.transform_expr(t.resolve_enum_shorthand(arg, enum_type))

	// Transform the receiver to apply smartcast if needed
	transformed_receiver := t.transform_expr(receiver)

	// Cast receiver to int: int(receiver)
	receiver_int := ast.CastExpr{
		typ:  ast.Ident{
			name: 'int'
		}
		expr: transformed_receiver
	}

	// Cast arg to int: int(flag)
	arg_int := ast.CastExpr{
		typ:  ast.Ident{
			name: 'int'
		}
		expr: resolved_arg
	}

	// receiver & flag
	and_expr := ast.InfixExpr{
		op:  .amp
		lhs: receiver_int
		rhs: arg_int
	}

	if method == 'has' {
		// (receiver & flag) != 0
		paren_pos := t.next_synth_pos()
		if int_obj := t.scope.lookup_parent('int', 0) {
			t.register_synth_type(paren_pos, int_obj.typ())
		}
		return ast.InfixExpr{
			op:  .ne
			lhs: ast.ParenExpr{
				expr: and_expr
				pos:  paren_pos
			}
			rhs: ast.BasicLiteral{
				kind:  .number
				value: '0'
			}
		}
	} else { // all
		// (receiver & flags) == int(flags)
		arg_int2 := ast.CastExpr{
			typ:  ast.Ident{
				name: 'int'
			}
			expr: resolved_arg
		}
		paren_pos := t.next_synth_pos()
		if int_obj := t.scope.lookup_parent('int', 0) {
			t.register_synth_type(paren_pos, int_obj.typ())
		}
		return ast.InfixExpr{
			op:  .eq
			lhs: ast.ParenExpr{
				expr: and_expr
				pos:  paren_pos
			}
			rhs: arg_int2
		}
	}
}

// try_transform_flag_enum_set_clear handles flag enum .set() and .clear() calls
// at the statement level, transforming them into compound assignment statements:
//   receiver.set(flag)   → receiver |= flag
//   receiver.clear(flag) → receiver &= ~flag
fn (mut t Transformer) try_transform_flag_enum_set_clear(stmt ast.ExprStmt) ?ast.Stmt {
	// Handle direct method call form: receiver.set(flag) / receiver.clear(flag)
	if stmt.expr is ast.CallExpr {
		call := stmt.expr as ast.CallExpr
		if call.lhs is ast.SelectorExpr {
			sel := call.lhs as ast.SelectorExpr
			method_name := sel.rhs.name
			if method_name in ['set', 'clear'] && call.args.len == 1 {
				receiver_type := t.get_enum_type(sel.lhs)
				if t.is_flag_enum_receiver(sel.lhs, receiver_type) {
					return t.make_flag_enum_assign(sel.lhs, method_name, call.args[0],
						receiver_type)
				}
			}
		}
		// Handle already-lowered form: Type__set(receiver, flag) / Type__clear(receiver, flag)
		if call.lhs is ast.Ident && call.args.len == 2 {
			name := call.lhs.name
			if name.ends_with('__set') || name.ends_with('__clear') {
				receiver_type := t.get_enum_type(call.args[0])
				if t.is_flag_enum_receiver(call.args[0], receiver_type) {
					method := if name.ends_with('__set') { 'set' } else { 'clear' }
					return t.make_flag_enum_assign(call.args[0], method, call.args[1],
						receiver_type)
				}
			}
		}
	}
	// Handle CallOrCastExpr form (single-arg method calls may be parsed this way)
	if stmt.expr is ast.CallOrCastExpr {
		coce := stmt.expr as ast.CallOrCastExpr
		if coce.lhs is ast.SelectorExpr {
			sel := coce.lhs as ast.SelectorExpr
			method_name := sel.rhs.name
			if method_name in ['set', 'clear'] {
				receiver_type := t.get_enum_type(sel.lhs)
				if t.is_flag_enum_receiver(sel.lhs, receiver_type) {
					return t.make_flag_enum_assign(sel.lhs, method_name, coce.expr, receiver_type)
				}
			}
		}
	}
	return none
}

// make_flag_enum_assign creates an AssignStmt for flag enum set/clear:
//   set:   receiver |= flag
//   clear: receiver &= ~flag
fn (mut t Transformer) make_flag_enum_assign(receiver ast.Expr, method string, arg ast.Expr, enum_type string) ast.Stmt {
	resolved_arg := t.resolve_enum_shorthand(arg, enum_type)
	transformed_receiver := t.transform_expr(receiver)
	transformed_arg := t.transform_expr(resolved_arg)

	if method == 'set' {
		// receiver |= flag
		return ast.AssignStmt{
			op:  .or_assign
			lhs: [ast.Expr(transformed_receiver)]
			rhs: [ast.Expr(transformed_arg)]
		}
	} else {
		// receiver &= ~flag
		return ast.AssignStmt{
			op:  .and_assign
			lhs: [ast.Expr(transformed_receiver)]
			rhs: [
				ast.Expr(ast.PrefixExpr{
					op:   .bit_not
					expr: transformed_arg
				}),
			]
		}
	}
}

// resolve_enum_shorthand resolves .member → EnumType.member
fn (t &Transformer) resolve_enum_shorthand(expr ast.Expr, enum_type string) ast.Expr {
	if expr is ast.SelectorExpr {
		sel := expr as ast.SelectorExpr
		// Check if it's a shorthand: .member (lhs is EmptyExpr or missing)
		if sel.lhs is ast.EmptyExpr {
			// Resolve to EnumType__member as an Ident (C-mangled name)
			return ast.Ident{
				name: '${enum_type}__${sel.rhs.name}'
				pos:  sel.pos
			}
		}
	}
	// For complex expressions (like flag1 | flag2), transform recursively
	if expr is ast.InfixExpr {
		infix := expr as ast.InfixExpr
		return ast.InfixExpr{
			op:  infix.op
			lhs: t.resolve_enum_shorthand(infix.lhs, enum_type)
			rhs: t.resolve_enum_shorthand(infix.rhs, enum_type)
			pos: infix.pos
		}
	}
	if expr is ast.ParenExpr {
		paren := expr as ast.ParenExpr
		return ast.ParenExpr{
			expr: t.resolve_enum_shorthand(paren.expr, enum_type)
			pos:  paren.pos
		}
	}
	return expr
}

// transform_array_with_enum_context transforms an array init, resolving enum shorthand using the given enum type
fn (mut t Transformer) transform_array_with_enum_context(arr ast.ArrayInitExpr, enum_type string) ast.Expr {
	mut exprs := []ast.Expr{cap: arr.exprs.len}
	for e in arr.exprs {
		// Resolve enum shorthand before transforming
		resolved := t.resolve_enum_shorthand(e, enum_type)
		exprs << t.transform_expr(resolved)
	}
	// Now create the transformed array init
	return t.transform_array_init_with_exprs(arr, exprs)
}

// transform_array_init_with_exprs transforms an array init using already-transformed expressions
fn (mut t Transformer) transform_array_init_with_exprs(arr ast.ArrayInitExpr, exprs []ast.Expr) ast.Expr {
	// Check if this is a fixed-size array
	mut is_fixed := false
	mut elem_type_expr := ast.empty_expr
	match arr.typ {
		ast.Type {
			if arr.typ is ast.ArrayFixedType {
				is_fixed = true
			} else if arr.typ is ast.ArrayType {
				elem_type_expr = arr.typ.elem_type
			}
		}
		else {}
	}
	// Also check for [x, y, z]! syntax - parser marks this with len: PostfixExpr{op: .not}
	if arr.len is ast.PostfixExpr {
		postfix := arr.len as ast.PostfixExpr
		if postfix.op == .not && postfix.expr is ast.EmptyExpr {
			is_fixed = true
		}
	}

	if is_fixed {
		return ast.ArrayInitExpr{
			typ:   arr.typ
			exprs: exprs
			init:  t.transform_expr(arr.init)
			cap:   arr.cap
			len:   arr.len
			pos:   arr.pos
		}
	}

	// Dynamic array: transform to builtin__new_array_from_c_array_noscan
	arr_len := exprs.len
	mut elem_type_name := 'int'
	mut elem_type_expr2 := elem_type_expr
	if elem_type_expr2 is ast.EmptyExpr && exprs.len > 0 {
		if arr_type := t.env.get_expr_type(arr.pos.id) {
			if arr_type is types.Array {
				tn := t.type_to_c_name(arr_type.elem_type)
				if tn != '' {
					elem_type_name = tn
					elem_type_expr2 = ast.Expr(ast.Ident{
						name: tn
					})
				}
			}
		}
		// If env lookup failed, try getting element type from the ORIGINAL first expression
		if elem_type_expr2 is ast.EmptyExpr && arr.exprs.len > 0 {
			if elem_type := t.get_expr_type(arr.exprs[0]) {
				tn := t.type_to_c_name(elem_type)
				if tn != '' {
					elem_type_name = tn
					elem_type_expr2 = ast.Expr(ast.Ident{
						name: tn
					})
				}
			}
		}
	}
	sizeof_arg := if elem_type_expr2 !is ast.EmptyExpr {
		elem_type_name = t.expr_to_type_name(elem_type_expr2)
		elem_type_expr2
	} else if exprs.len > 0 {
		first := exprs[0]
		if first is ast.BasicLiteral {
			if first.kind == .number {
				if first.value.contains('.') || first.value.contains('e')
					|| first.value.contains('E') {
					elem_type_name = 'f64'
				} else {
					elem_type_name = 'int'
				}
			} else if first.kind == .string {
				elem_type_name = 'string'
			}
			ast.Expr(ast.Ident{
				name: elem_type_name
			})
		} else if first is ast.StringLiteral {
			elem_type_name = 'string'
			ast.Expr(ast.Ident{
				name: 'string'
			})
		} else if first is ast.SelectorExpr {
			// For qualified enum values, use int for sizeof
			elem_type_name = 'int'
			ast.Expr(ast.Ident{
				name: 'int'
			})
		} else if first is ast.InitExpr {
			// Struct literal - get the type name from the struct type
			init_type_name := t.expr_to_type_name(first.typ)
			if init_type_name != '' {
				elem_type_name = init_type_name
				ast.Expr(ast.Ident{
					name: init_type_name
				})
			} else {
				exprs[0]
			}
		} else {
			exprs[0]
		}
	} else {
		ast.Expr(ast.Ident{
			name: 'int'
		})
	}

	// Create proper array type for the inner ArrayInitExpr
	inner_array_typ := ast.Type(ast.ArrayType{
		elem_type: ast.Ident{
			name: elem_type_name
		}
	})

	return ast.CallExpr{
		lhs:  ast.Ident{
			name: 'builtin__new_array_from_c_array_noscan'
		}
		args: [
			ast.Expr(ast.BasicLiteral{
				kind:  .number
				value: '${arr_len}'
			}),
			ast.Expr(ast.BasicLiteral{
				kind:  .number
				value: '${arr_len}'
			}),
			ast.Expr(ast.KeywordOperator{
				op:    .key_sizeof
				exprs: [sizeof_arg]
			}),
			ast.Expr(ast.ArrayInitExpr{
				typ:   ast.Expr(inner_array_typ)
				exprs: exprs
			}),
		]
		pos:  arr.pos
	}
}

// rename_substr_to_checked renames a string__substr call to string__substr_with_check.
// Used for string range with or-blocks: s[0..20] or { 'fallback' } needs the checked
// variant which returns !string (Result) instead of plain string.
fn (t &Transformer) rename_substr_to_checked(expr ast.Expr) ast.Expr {
	if expr is ast.CallExpr {
		if expr.lhs is ast.Ident && expr.lhs.name == 'string__substr' {
			return ast.CallExpr{
				lhs:  ast.Ident{
					name: 'string__substr_with_check'
				}
				args: expr.args
			}
		}
	}
	return expr
}

// is_string_expr returns true if the expression is known to be a string
fn (t &Transformer) is_string_expr(expr ast.Expr) bool {
	if expr is ast.StringLiteral {
		// Check for c-strings which are char*, not string
		return !expr.value.starts_with("c'")
	}
	if expr is ast.StringInterLiteral {
		return true
	}
	if expr is ast.BasicLiteral {
		return expr.kind == .string
	}
	if expr is ast.ComptimeExpr {
		// Compile-time expressions like @FN, @FILE, @MOD evaluate to strings
		if expr.expr is ast.Ident {
			name := (expr.expr as ast.Ident).name
			return name in ['FN', 'FILE', 'MOD', 'STRUCT', 'METHOD', 'LOCATION', 'FUNCTION']
		}
	}
	if expr is ast.CastExpr {
		// Check if casting to string type
		if expr.typ is ast.Ident {
			return expr.typ.name == 'string'
		}
	}
	if expr is ast.Ident {
		// Check for comptime string identifiers like @FN, @FILE, @MOD
		if expr.name.starts_with('@') {
			return expr.name in ['@FN', '@FILE', '@MOD', '@STRUCT', '@METHOD', '@LOCATION',
				'@FUNCTION', '@VMODROOT']
		}
		// Check if variable type is string via scope lookup
		var_type_name := t.get_var_type_name(expr.name)
		if var_type_name == 'string' {
			return true
		}
		// Use type environment to look up the identifier's type
		if mut scope := t.get_current_scope() {
			if obj := scope.lookup_parent(expr.name, 0) {
				typ := obj.typ()
				if typ is types.String {
					return true
				}
				// Also check for struct named 'string' (V's string type)
				if typ is types.Struct && (typ as types.Struct).name == 'string' {
					return true
				}
			}
		}
	}
	if expr is ast.ParenExpr {
		return t.is_string_expr(expr.expr)
	}
	if expr is ast.SelectorExpr {
		// Check for module-qualified constants (e.g., os.path_separator)
		if expr.lhs is ast.Ident {
			mod_name := (expr.lhs as ast.Ident).name
			const_name := expr.rhs.name
			// Try to look up the constant in the module's scope
			if mut mod_scope := t.get_module_scope(mod_name) {
				if obj := mod_scope.lookup_parent(const_name, 0) {
					typ := obj.typ()
					if typ is types.String {
						return true
					}
					if typ is types.Struct && (typ as types.Struct).name == 'string' {
						return true
					}
				}
			}
		}
		// Try to look up the type of the field using the environment
		if lhs_type := t.get_expr_type(expr.lhs) {
			base_type := if lhs_type is types.Pointer {
				lhs_type.base_type
			} else {
				lhs_type
			}
			if base_type is types.Struct {
				for field in base_type.fields {
					if field.name == expr.rhs.name {
						if field.typ is types.String {
							return true
						}
						if field.typ is types.Struct {
							field_struct := field.typ as types.Struct
							if field_struct.name == 'string' {
								return true
							}
						}
					}
				}
			}
		}
		// Fallback: Check field names that are typically strings
		// Only use this for common string field names
		if expr.rhs.name in ['name', 'str', 'msg'] {
			return true
		}
	}
	if expr is ast.UnsafeExpr {
		// Check the last statement's expression inside unsafe blocks
		// e.g., unsafe { s.substr_unsafe(i, j) }
		if expr.stmts.len > 0 {
			last_stmt := expr.stmts[expr.stmts.len - 1]
			if last_stmt is ast.ExprStmt {
				return t.is_string_expr(last_stmt.expr)
			}
		}
	}
	if expr is ast.IndexExpr {
		// String slicing: s[a..b] returns string if s is string
		if expr.expr is ast.RangeExpr {
			return t.is_string_expr(expr.lhs)
		}
		// Array indexing: arr[i] where arr is []string returns string
		if expr.lhs is ast.Ident {
			arr_name := (expr.lhs as ast.Ident).name
			arr_type := t.get_var_type_name(arr_name)
			if arr_type == 'Array_string' {
				return true
			}
		}
		// Use get_expr_type which handles IndexExpr and returns the element type
		if elem_type := t.get_expr_type(expr) {
			if elem_type is types.String {
				return true
			}
			if elem_type is types.Struct && (elem_type as types.Struct).name == 'string' {
				return true
			}
		}
	}
	if expr is ast.InfixExpr {
		// For + on strings, result is string
		if expr.op == .plus && t.is_string_expr(expr.lhs) {
			return true
		}
	}
	if expr is ast.CallExpr {
		// Check method calls that return string using types.Environment
		if expr.lhs is ast.SelectorExpr {
			sel := expr.lhs as ast.SelectorExpr
			method_name := sel.rhs.name
			// First check for module-qualified function calls (e.g., os.user_os())
			// If LHS is an Ident, it could be a module name
			if sel.lhs is ast.Ident {
				mod_name := (sel.lhs as ast.Ident).name
				// Try looking up as a module-qualified function
				if fn_type := t.env.lookup_fn(mod_name, method_name) {
					if return_type := fn_type.get_return_type() {
						if return_type is types.String {
							return true
						}
						if return_type is types.Struct
							&& (return_type as types.Struct).name == 'string' {
							return true
						}
					}
				}
			}
			// Try method lookup
			if receiver_type := t.get_expr_type(sel.lhs) {
				type_name := t.get_type_name(receiver_type)
				if fn_type := t.env.lookup_method(type_name, method_name) {
					if return_type := fn_type.get_return_type() {
						if return_type is types.String {
							return true
						}
						if return_type is types.Struct
							&& (return_type as types.Struct).name == 'string' {
							return true
						}
					}
				}
			}
			// Check for array methods that return element type (pop, first, last)
			// If receiver is []string, these methods return string
			if method_name in ['pop', 'first', 'last'] {
				if sel.lhs is ast.Ident {
					receiver_name := (sel.lhs as ast.Ident).name
					receiver_type := t.get_var_type_name(receiver_name)
					if receiver_type == 'Array_string' {
						return true
					}
				}
			}
			// Fallback: check known string-returning methods
			if t.is_string_returning_method(method_name) {
				return true
			}
			// Also check if receiver is string and method typically returns string
			if t.is_string_expr(sel.lhs) && method_name in ['clone', 'str', 'string'] {
				return true
			}
		}
		// Check function return type using environment
		if expr.lhs is ast.Ident {
			fn_name := expr.lhs.name
			// Check for already-transformed string functions
			if fn_name.starts_with('string__') && fn_name !in ['string__bytes', 'string__vbytes'] {
				// string__ prefix functions return string (string__plus, string__repeat, etc.)
				// except string__bytes/string__vbytes which return []u8
				return true
			}
			// Try to find the function in the current module's scope
			if mut scope := t.get_current_scope() {
				if obj := scope.lookup_parent(fn_name, 0) {
					typ := obj.typ()
					if typ is types.FnType {
						if return_type := typ.get_return_type() {
							if return_type is types.String {
								return true
							}
							if return_type is types.Struct
								&& (return_type as types.Struct).name == 'string' {
								return true
							}
						}
					}
				}
			}
			// Fallback: check if function name is known to return string
			if t.is_string_returning_fn(fn_name) {
				return true
			}
			// Handle cross-module function calls like os__user_os()
			// Parse module prefix (e.g., os__user_os -> module: os, fn: user_os)
			if fn_name.contains('__') {
				parts := fn_name.split('__')
				if parts.len >= 2 {
					mod_name := parts[0]
					actual_fn := parts[1..].join('__')
					// Use environment's lookup_fn which checks the module's scope
					if fn_type := t.env.lookup_fn(mod_name, actual_fn) {
						if return_type := fn_type.get_return_type() {
							if return_type is types.String {
								return true
							}
							if return_type is types.Struct
								&& (return_type as types.Struct).name == 'string' {
								return true
							}
						}
					}
					// Fallback: check if function name is known to return string
					if t.is_string_returning_fn(actual_fn) {
						return true
					}
				}
			}
		}
	}
	if expr is ast.CallOrCastExpr {
		// Check method calls for CallOrCastExpr (single-arg method calls like 'foo'.repeat(5))
		if expr.lhs is ast.SelectorExpr {
			sel := expr.lhs as ast.SelectorExpr
			method_name := sel.rhs.name
			// First check for module-qualified function calls (e.g., os.user_os())
			if sel.lhs is ast.Ident {
				mod_name := (sel.lhs as ast.Ident).name
				if fn_type := t.env.lookup_fn(mod_name, method_name) {
					if return_type := fn_type.get_return_type() {
						if return_type is types.String {
							return true
						}
						if return_type is types.Struct
							&& (return_type as types.Struct).name == 'string' {
							return true
						}
					}
				}
			}
			// Try method lookup
			if receiver_type := t.get_expr_type(sel.lhs) {
				type_name := t.get_type_name(receiver_type)
				if fn_type := t.env.lookup_method(type_name, method_name) {
					if return_type := fn_type.get_return_type() {
						if return_type is types.String {
							return true
						}
						if return_type is types.Struct
							&& (return_type as types.Struct).name == 'string' {
							return true
						}
					}
				}
			}
			// Fallback: check known string-returning methods
			if t.is_string_returning_method(method_name) {
				return true
			}
			// Also check if receiver is string and method typically returns string
			if t.is_string_expr(sel.lhs) && method_name in ['clone', 'str', 'string'] {
				return true
			}
		}
		// Check function return type for CallOrCastExpr (single-arg calls)
		if expr.lhs is ast.Ident {
			fn_name := expr.lhs.name
			// Check for already-transformed string functions
			if fn_name.starts_with('string__') {
				return true
			}
			if mut scope := t.get_current_scope() {
				if obj := scope.lookup_parent(fn_name, 0) {
					typ := obj.typ()
					if typ is types.FnType {
						if return_type := typ.get_return_type() {
							if return_type is types.String {
								return true
							}
							if return_type is types.Struct
								&& (return_type as types.Struct).name == 'string' {
								return true
							}
						}
					}
				}
			}
			// Fallback: check if function name is known to return string
			if t.is_string_returning_fn(fn_name) {
				return true
			}
			// Handle cross-module function calls like os__user_os()
			if fn_name.contains('__') {
				parts := fn_name.split('__')
				if parts.len >= 2 {
					mod_name := parts[0]
					actual_fn := parts[1..].join('__')
					if fn_type := t.env.lookup_fn(mod_name, actual_fn) {
						if return_type := fn_type.get_return_type() {
							if return_type is types.String {
								return true
							}
							if return_type is types.Struct
								&& (return_type as types.Struct).name == 'string' {
								return true
							}
						}
					}
					// Fallback: check if function name is known to return string
					if t.is_string_returning_fn(actual_fn) {
						return true
					}
				}
			}
		}
	}
	if expr is ast.IfExpr {
		// For ternary if-expressions, check if both branches are strings
		// Check 'then' branch (stmts - last stmt should be an expression)
		if expr.stmts.len > 0 {
			last_stmt := expr.stmts[expr.stmts.len - 1]
			if last_stmt is ast.ExprStmt {
				// Use context-aware check that looks at assignments within this block
				if !t.is_string_expr_in_block(last_stmt.expr, expr.stmts) {
					return false
				}
			}
		}
		// Check 'else' branch
		if expr.else_expr is ast.IfExpr {
			if !t.is_string_expr(expr.else_expr) {
				return false
			}
		} else if expr.else_expr !is ast.EmptyExpr {
			// else_expr could be a single expression
			if !t.is_string_expr(expr.else_expr) {
				return false
			}
		}
		// If we get here and had at least one branch, treat as string
		return expr.stmts.len > 0
	}
	// Fallback: use type environment for any expression type
	if elem_type := t.get_expr_type(expr) {
		if elem_type is types.String {
			return true
		}
		if elem_type is types.Struct && (elem_type as types.Struct).name == 'string' {
			return true
		}
	}
	return false
}

// is_string_expr_in_block checks if an expression is a string, with context from block statements
fn (t &Transformer) is_string_expr_in_block(expr ast.Expr, stmts []ast.Stmt) bool {
	// Handle IndexExpr into local array variables within this block
	if expr is ast.IndexExpr {
		if expr.lhs is ast.Ident {
			arr_name := (expr.lhs as ast.Ident).name
			arr_type := t.find_var_type_in_stmts(stmts, arr_name)
			if arr_type == 'Array_string' {
				return true
			}
		}
	}
	// Fall back to regular is_string_expr
	return t.is_string_expr(expr)
}

// is_string_returning_fn returns true if a function is known to return a string
fn (t &Transformer) is_string_returning_fn(fn_name string) bool {
	// Known string-returning functions
	if fn_name in ['string__plus', 'string__plus_two', 'string__substr', 'string__substr_unsafe',
		'string__repeat'] {
		return true
	}
	// String module functions generally return strings (except bytes/vbytes which return []u8)
	if fn_name.starts_with('string__') && fn_name !in ['string__bytes', 'string__vbytes'] {
		return true
	}
	// Check function return type using scope lookup
	if ret_type := t.get_fn_return_type(fn_name) {
		if ret_type.name() == 'string' {
			return true
		}
	}
	// Recognize functions by naming pattern
	if fn_name.ends_with('_to_string') || fn_name.ends_with('__str') {
		return true
	}
	// int/u8/etc hex() method gets converted to int__hex etc
	if fn_name.ends_with('__hex') || fn_name.ends_with('__str') {
		return true
	}
	return false
}

// is_string_returning_method returns true if a method is known to return a string
fn (t &Transformer) is_string_returning_method(method_name string) bool {
	// Common string methods that return string
	return method_name in [
		'str',
		'string',
		'to_upper',
		'to_lower',
		'capitalize',
		'uncapitalize',
		'trim',
		'trim_left',
		'trim_right',
		'trim_space',
		'strip_margin',
		'replace',
		'replace_once',
		'substr',
		'substr_unsafe',
		'repeat',
		'reverse',
		'after',
		'before',
		'all_before',
		'all_after',
		'all_before_last',
		'all_after_last',
		'join',
		'ascii_str',
		'hex',
		'clone',
		'bytestr',
		// Code generation methods that return string
		'gen',
		'name',
		// Error message methods
		'posix_get_error_msg',
		'get_error_msg',
	]
}

// get_str_fn_name_for_expr returns the str function name for an expression's type.
// For example: []int -> Array_int_str, map[string]int -> Map_string_int_str
fn (t &Transformer) get_str_fn_name_for_expr(expr ast.Expr) ?string {
	// First try to infer array type
	if array_type := t.get_array_type_str(expr) {
		// array_type is like 'Array_int', so append '_str'
		return '${array_type}_str'
	}
	// Try to infer map type
	if map_type := t.get_map_type_for_expr(expr) {
		// map_type is like 'Map_string_int', so append '_str'
		return '${map_type}_str'
	}
	// Try to get type from expression
	if typ := t.get_expr_type(expr) {
		return t.get_str_fn_name_for_type(typ)
	}
	// Handle ArrayInitExpr directly for inline array literals
	if expr is ast.ArrayInitExpr {
		// Get element type from first element or type annotation
		elem_type := t.get_array_init_elem_type(expr)
		if elem_type != '' {
			return 'Array_${elem_type}_str'
		}
		return 'Array_int_str' // Default fallback
	}
	return none
}

// StrFnInfo holds information about an auto-generated str function
struct StrFnInfo {
	str_fn_name string
	elem_type   string
}

// get_str_fn_info_for_expr returns the str function name and element type info for auto-generation.
// Returns StrFnInfo with str_fn_name and elem_type where elem_type is the element type for arrays.
fn (mut t Transformer) get_str_fn_info_for_expr(expr ast.Expr) StrFnInfo {
	// First try to infer array type
	if array_type := t.get_array_type_str(expr) {
		// array_type is like 'Array_int'
		elem_type := array_type['Array_'.len..]
		return StrFnInfo{
			str_fn_name: '${array_type}_str'
			elem_type:   elem_type
		}
	}
	// Try to infer map type
	if map_type := t.get_map_type_for_expr(expr) {
		// map_type is like 'Map_string_int'
		return StrFnInfo{
			str_fn_name: '${map_type}_str'
			elem_type:   map_type
		}
	}
	// Handle ArrayInitExpr directly for inline array literals
	if expr is ast.ArrayInitExpr {
		elem_type := t.get_array_init_elem_type(expr)
		if elem_type != '' {
			return StrFnInfo{
				str_fn_name: 'Array_${elem_type}_str'
				elem_type:   elem_type
			}
		}
		return StrFnInfo{
			str_fn_name: 'Array_int_str'
			elem_type:   'int'
		}
	}
	// Handle enum, struct, and primitive types via type lookup
	if typ := t.get_expr_type(expr) {
		if str_fn_name := t.get_str_fn_name_for_type(typ) {
			return StrFnInfo{
				str_fn_name: str_fn_name
				elem_type:   typ.name()
			}
		}
	}
	return StrFnInfo{}
}

// generate_str_functions generates FnDecl AST nodes for needed auto str functions.
// For arrays: generates a function that iterates over elements and calls their str methods.
fn (mut t Transformer) generate_str_functions() []ast.Stmt {
	mut result := []ast.Stmt{cap: t.needed_str_fns.len}
	for fn_name, elem_type in t.needed_str_fns {
		// Generate array str function (skip fixed arrays - they need different handling)
		if fn_name.starts_with('Array_') && !fn_name.starts_with('Array_fixed_') {
			result << t.generate_array_str_fn(fn_name, elem_type)
		}
	}
	return result
}

enum ArrayMethodKind {
	contains
	index
	last_index
}

fn (mut t Transformer) generate_array_method_functions() []ast.Stmt {
	mut result := []ast.Stmt{cap: t.needed_array_contains_fns.len + t.needed_array_index_fns.len +
		t.needed_array_last_index_fns.len}
	mut contains_names := t.needed_array_contains_fns.keys()
	contains_names.sort()
	for fn_name in contains_names {
		result << t.generate_array_method_fn(fn_name, t.needed_array_contains_fns[fn_name],
			.contains)
	}
	mut index_names := t.needed_array_index_fns.keys()
	index_names.sort()
	for fn_name in index_names {
		result << t.generate_array_method_fn(fn_name, t.needed_array_index_fns[fn_name],
			.index)
	}
	mut last_index_names := t.needed_array_last_index_fns.keys()
	last_index_names.sort()
	for fn_name in last_index_names {
		result << t.generate_array_method_fn(fn_name, t.needed_array_last_index_fns[fn_name],
			.last_index)
	}
	return result
}

fn (mut t Transformer) generate_array_method_len_expr(info ArrayMethodInfo) ast.Expr {
	if info.is_fixed {
		return ast.Expr(ast.BasicLiteral{
			kind:  .number
			value: info.fixed_len.str()
		})
	}
	return t.synth_selector(ast.Ident{ name: 'a' }, 'len', types.Type(types.int_))
}

fn (mut t Transformer) generate_array_method_elem_expr(info ArrayMethodInfo, idx_expr ast.Expr) ast.Expr {
	if info.is_fixed {
		return ast.Expr(ast.IndexExpr{
			lhs:  ast.Ident{
				name: 'a'
			}
			expr: idx_expr
		})
	}
	return ast.Expr(ast.PrefixExpr{
		op:   .mul
		expr: ast.CastExpr{
			typ:  ast.PrefixExpr{
				op:   .amp
				expr: ast.Ident{
					name: info.elem_type
				}
			}
			expr: ast.CallExpr{
				lhs:  ast.Ident{
					name: 'array__get'
				}
				args: [
					ast.Expr(ast.Ident{
						name: 'a'
					}),
					idx_expr,
				]
			}
		}
	})
}

fn (mut t Transformer) generate_array_method_match_expr(info ArrayMethodInfo, idx_expr ast.Expr) ast.Expr {
	elem_expr := t.generate_array_method_elem_expr(info, idx_expr)
	if info.elem_type == 'string' {
		return ast.Expr(ast.CallExpr{
			lhs:  ast.Ident{
				name: 'string__eq'
			}
			args: [
				elem_expr,
				ast.Expr(ast.Ident{
					name: 'v'
				}),
			]
		})
	}
	if info.elem_type.starts_with('Array_') {
		return ast.Expr(ast.CallExpr{
			lhs:  ast.Ident{
				name: 'array__eq'
			}
			args: [
				ast.Expr(ast.ParenExpr{
					expr: elem_expr
				}),
				ast.Expr(ast.Ident{
					name: 'v'
				}),
			]
		})
	}
	return ast.Expr(ast.InfixExpr{
		op:  .eq
		lhs: elem_expr
		rhs: ast.Ident{
			name: 'v'
		}
	})
}

fn (mut t Transformer) generate_array_method_loop_stmt(info ArrayMethodInfo, kind ArrayMethodKind, loop_body []ast.Stmt) ast.Stmt {
	mut init_rhs := ast.Expr(ast.BasicLiteral{
		kind:  .number
		value: '0'
	})
	mut cond_op := token.Token.lt
	mut cond_rhs := t.generate_array_method_len_expr(info)
	mut post_op := token.Token.plus_assign
	mut post_rhs := ast.Expr(ast.BasicLiteral{
		kind:  .number
		value: '1'
	})
	if kind == .last_index {
		init_rhs = if info.is_fixed {
			ast.Expr(ast.BasicLiteral{
				kind:  .number
				value: (info.fixed_len - 1).str()
			})
		} else {
			ast.Expr(ast.InfixExpr{
				op:  .minus
				lhs: t.synth_selector(ast.Ident{ name: 'a' }, 'len', types.Type(types.int_))
				rhs: ast.BasicLiteral{
					kind:  .number
					value: '1'
				}
			})
		}
		cond_op = .ge
		cond_rhs = ast.Expr(ast.BasicLiteral{
			kind:  .number
			value: '0'
		})
		post_op = .minus_assign
	}
	return ast.Stmt(ast.ForStmt{
		init:  ast.AssignStmt{
			op:  .decl_assign
			lhs: [
				ast.Expr(ast.Ident{
					name: 'i'
				}),
			]
			rhs: [init_rhs]
		}
		cond:  ast.InfixExpr{
			op:  cond_op
			lhs: ast.Ident{
				name: 'i'
			}
			rhs: cond_rhs
		}
		post:  ast.AssignStmt{
			op:  post_op
			lhs: [
				ast.Expr(ast.Ident{
					name: 'i'
				}),
			]
			rhs: [post_rhs]
		}
		stmts: loop_body
	})
}

fn (mut t Transformer) generate_array_method_fn(fn_name string, info ArrayMethodInfo, kind ArrayMethodKind) ast.Stmt {
	param_a := ast.Parameter{
		name: 'a'
		typ:  ast.Ident{
			name: info.array_type
		}
	}
	param_v := ast.Parameter{
		name: 'v'
		typ:  ast.Ident{
			name: info.elem_type
		}
	}
	// Register a function scope so cleanc can resolve parameter types via scope lookup.
	t.register_generated_fn_scope(fn_name, 'builtin', [param_a, param_v])
	idx_expr := ast.Expr(ast.Ident{
		name: 'i'
	})
	cond_expr := t.generate_array_method_match_expr(info, idx_expr)
	match_ret := if kind == .contains {
		ast.Expr(ast.Keyword{
			tok: .key_true
		})
	} else {
		idx_expr
	}
	mut loop_body := []ast.Stmt{}
	loop_body << ast.ExprStmt{
		expr: ast.IfExpr{
			cond:  cond_expr
			stmts: [
				ast.Stmt(ast.ReturnStmt{
					exprs: [match_ret]
				}),
			]
		}
	}
	mut body_stmts := []ast.Stmt{}
	body_stmts << t.generate_array_method_loop_stmt(info, kind, loop_body)
	fallback_ret := if kind == .contains {
		ast.Expr(ast.Keyword{
			tok: .key_false
		})
	} else {
		ast.Expr(ast.BasicLiteral{
			kind:  .number
			value: '-1'
		})
	}
	body_stmts << ast.ReturnStmt{
		exprs: [fallback_ret]
	}
	return_type_name := if kind == .contains { 'bool' } else { 'int' }
	return ast.Stmt(ast.FnDecl{
		name:       fn_name
		is_public:  false
		is_method:  false
		is_static:  false
		attributes: []ast.Attribute{}
		typ:        ast.FnType{
			params:      [param_a, param_v]
			return_type: ast.Ident{
				name: return_type_name
			}
		}
		stmts:      body_stmts
	})
}

// generate_array_str_fn generates a str function for an array type.
// Example for Array_int_str:
//   fn Array_int_str(a Array_int) string {
//       mut sb := strings__new_builder(2 + a.len * 10)
//       strings__Builder__write_string(&sb, "[")
//       for i := 0; i < a.len; i++ {
//           if i > 0 { strings__Builder__write_string(&sb, ", ") }
//           strings__Builder__write_string(&sb, int_str(a.data[i]))
//       }
//       strings__Builder__write_string(&sb, "]")
//       return strings__Builder__str(&sb)
//   }
fn (mut t Transformer) generate_array_str_fn(fn_name string, elem_type string) ast.Stmt {
	// Create parameter: a Array_int
	array_type_name := fn_name[..fn_name.len - 4] // Remove '_str' suffix: 'Array_int_str' -> 'Array_int'
	param_a := ast.Parameter{
		name: 'a'
		typ:  ast.Ident{
			name: array_type_name
		}
	}
	// Register a function scope so cleanc can resolve parameter types via scope lookup.
	t.register_generated_fn_scope(fn_name, 'builtin', [param_a])

	// Get element str function name.
	// Auto-generated helper functions (Array_, Map_) use single underscore _str suffix.
	// Real type methods use double underscore __str suffix.
	// For pointer element types (e.g. Coordptr), strip 'ptr' suffix to get base type str fn.
	mut resolved_elem_type := elem_type
	if elem_type.ends_with('ptr') && elem_type != 'voidptr' && elem_type != 'charptr'
		&& elem_type != 'byteptr' {
		resolved_elem_type = elem_type[..elem_type.len - 3]
	}
	elem_str_fn := if resolved_elem_type.starts_with('Array_')
		|| resolved_elem_type.starts_with('Map_') {
		'${resolved_elem_type}_str'
	} else {
		'${resolved_elem_type}__str'
	}

	// Build the function body statements
	mut body_stmts := []ast.Stmt{}

	// mut sb := strings__new_builder(2 + a.len * 10)
	body_stmts << ast.AssignStmt{
		op:  .decl_assign
		lhs: [
			ast.Expr(ast.ModifierExpr{
				kind: .key_mut
				expr: ast.Ident{
					name: 'sb'
				}
			}),
		]
		rhs: [
			ast.Expr(ast.CallExpr{
				lhs:  ast.Ident{
					name: 'strings__new_builder'
				}
				args: [
					ast.Expr(ast.InfixExpr{
						op:  .plus
						lhs: ast.BasicLiteral{
							kind:  .number
							value: '2'
						}
						rhs: ast.InfixExpr{
							op:  .mul
							lhs: t.synth_selector(ast.Ident{ name: 'a' }, 'len', types.Type(types.int_))
							rhs: ast.BasicLiteral{
								kind:  .number
								value: '10'
							}
						}
					}),
				]
			}),
		]
	}

	// strings__Builder__write_string(&sb, "[")
	body_stmts << ast.ExprStmt{
		expr: ast.CallExpr{
			lhs:  ast.Ident{
				name: 'strings__Builder__write_string'
			}
			args: [
				ast.Expr(ast.PrefixExpr{
					op:   .amp
					expr: ast.Ident{
						name: 'sb'
					}
				}),
				ast.Expr(ast.StringLiteral{
					kind:  .v
					value: '['
				}),
			]
		}
	}

	// for i := 0; i < a.len; i++ { ... }
	// Build the for loop body
	mut for_body := []ast.Stmt{}

	// if i > 0 { strings__Builder__write_string(&sb, ", ") }
	for_body << ast.ExprStmt{
		expr: ast.IfExpr{
			cond:  ast.InfixExpr{
				op:  .gt
				lhs: ast.Ident{
					name: 'i'
				}
				rhs: ast.BasicLiteral{
					kind:  .number
					value: '0'
				}
			}
			stmts: [
				ast.Stmt(ast.ExprStmt{
					expr: ast.CallExpr{
						lhs:  ast.Ident{
							name: 'strings__Builder__write_string'
						}
						args: [
							ast.Expr(ast.PrefixExpr{
								op:   .amp
								expr: ast.Ident{
									name: 'sb'
								}
							}),
							ast.Expr(ast.StringLiteral{
								kind:  .v
								value: ', '
							}),
						]
					}
				}),
			]
		}
	}

	// strings__Builder__write_string(&sb, elem_str(*(elem_type*)array__get(a, i)))
	for_body << ast.ExprStmt{
		expr: ast.CallExpr{
			lhs:  ast.Ident{
				name: 'strings__Builder__write_string'
			}
			args: [
				ast.Expr(ast.PrefixExpr{
					op:   .amp
					expr: ast.Ident{
						name: 'sb'
					}
				}),
				// elem_str(*(elem_type*)array__get(a, i))
				ast.Expr(ast.CallExpr{
					lhs:  ast.Ident{
						name: elem_str_fn
					}
					args: [
						ast.Expr(ast.PrefixExpr{
							op:   .mul
							expr: ast.CastExpr{
								typ:  ast.PrefixExpr{
									op:   .amp
									expr: ast.Ident{
										name: elem_type
									}
								}
								expr: ast.CallExpr{
									lhs:  ast.Ident{
										name: 'array__get'
									}
									args: [
										ast.Expr(ast.Ident{
											name: 'a'
										}),
										ast.Expr(ast.Ident{
											name: 'i'
										}),
									]
								}
							}
						}),
					]
				}),
			]
		}
	}

	// for loop: for i := 0; i < a.len; i++ { ... }
	body_stmts << ast.ForStmt{
		init:  ast.AssignStmt{
			op:  .decl_assign
			lhs: [ast.Expr(ast.Ident{
				name: 'i'
			})]
			rhs: [ast.Expr(ast.BasicLiteral{
				kind:  .number
				value: '0'
			})]
		}
		cond:  ast.InfixExpr{
			op:  .lt
			lhs: ast.Ident{
				name: 'i'
			}
			rhs: t.synth_selector(ast.Ident{ name: 'a' }, 'len', types.Type(types.int_))
		}
		post:  ast.AssignStmt{
			op:  .plus_assign
			lhs: [ast.Expr(ast.Ident{
				name: 'i'
			})]
			rhs: [ast.Expr(ast.BasicLiteral{
				kind:  .number
				value: '1'
			})]
		}
		stmts: for_body
	}

	// strings__Builder__write_string(&sb, "]")
	body_stmts << ast.ExprStmt{
		expr: ast.CallExpr{
			lhs:  ast.Ident{
				name: 'strings__Builder__write_string'
			}
			args: [
				ast.Expr(ast.PrefixExpr{
					op:   .amp
					expr: ast.Ident{
						name: 'sb'
					}
				}),
				ast.Expr(ast.StringLiteral{
					kind:  .v
					value: ']'
				}),
			]
		}
	}

	// return strings__Builder__str(&sb)
	body_stmts << ast.ReturnStmt{
		exprs: [
			ast.Expr(ast.CallExpr{
				lhs:  ast.Ident{
					name: 'strings__Builder__str'
				}
				args: [
					ast.Expr(ast.PrefixExpr{
						op:   .amp
						expr: ast.Ident{
							name: 'sb'
						}
					}),
				]
			}),
		]
	}

	// Create the function declaration
	return ast.FnDecl{
		name:       fn_name
		is_public:  false
		is_method:  false
		is_static:  false
		attributes: []ast.Attribute{}
		typ:        ast.FnType{
			params:      [param_a]
			return_type: ast.Ident{
				name: 'string'
			}
		}
		stmts:      body_stmts
	}
}
