module main

fn main() {
	fa := get_fn_a()
	fb := get_fn_b()
	println(fa())
	println(fb())
}
